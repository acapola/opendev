﻿/*
Hamming code EDC/ECC modules library
*/
/////////////////////////////////////////////////////////////////////////////////////////////////
// *_min_width modules: use the least possible EDC bits
/////////////////////////////////////////////////////////////////////////////////////////////////
module edc_hc_4_min_width (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [3-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [3-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_7_4_f
//Compute 3 bits Error Detection Code from a 4 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 16 valid code words out of 128 therefore 87% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: xx x (3 inputs)
//  syndrom[1]: x xx (3 inputs)
//  syndrom[2]:  xxx (3 inputs)
//Input usage report:
//  input bit 0 used 2 times (syndrom bits 0 1)
//  input bit 1 used 2 times (syndrom bits 0 2)
//  input bit 2 used 2 times (syndrom bits 1 2)
//  input bit 3 used 3 times (syndrom bits 0 1 2)
function [3-1:0] hamming_code_7_4_f;
    input [4-1:0] in;
    reg [3-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[3];//3 inputs
        syndrom[1] = in[0]^in[2]^in[3];//3 inputs
        syndrom[2] = in[1]^in[2]^in[3];//3 inputs
        hamming_code_7_4_f = syndrom;
    end
endfunction
wire [3-1:0] stored_data_edc = hamming_code_7_4_f(i_stored_data);
wire [3-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_4_min_width (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: xxx  (3 inputs)
//  syndrom[1]: xx x (3 inputs)
//  syndrom[2]: x xx (3 inputs)
//  syndrom[3]:  xxx (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 1 3)
//  input bit 2 used 3 times (syndrom bits 0 2 3)
//  input bit 3 used 3 times (syndrom bits 1 2 3)
function [4-1:0] extended_hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[2];//3 inputs
        syndrom[1] = in[0]^in[1]^in[3];//3 inputs
        syndrom[2] = in[0]^in[2]^in[3];//3 inputs
        syndrom[3] = in[1]^in[2]^in[3];//3 inputs
        extended_hamming_code_8_4_f = syndrom;
    end
endfunction
wire [4-1:0] stored_data_edc = extended_hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_4_min_width (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [4-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: xxx  (3 inputs)
//  syndrom[1]: xx x (3 inputs)
//  syndrom[2]: x xx (3 inputs)
//  syndrom[3]:  xxx (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 1 3)
//  input bit 2 used 3 times (syndrom bits 0 2 3)
//  input bit 3 used 3 times (syndrom bits 1 2 3)
function [4-1:0] extended_hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[2];//3 inputs
        syndrom[1] = in[0]^in[1]^in[3];//3 inputs
        syndrom[2] = in[0]^in[2]^in[3];//3 inputs
        syndrom[3] = in[1]^in[2]^in[3];//3 inputs
        extended_hamming_code_8_4_f = syndrom;
    end
endfunction
function [2+4-1:0] extended_hamming_code_8_4_f_correction_pattern_f;
    input [4-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [4-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {4{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			4'b0000: begin
				correctable_error = 1'b0;
				correction_pattern = {4{1'b0}};
			end	
			4'b0111: begin
				correction_pattern = {4{1'b0}};correction_pattern[0]=1'b1;
			end
			4'b1011: begin
				correction_pattern = {4{1'b0}};correction_pattern[1]=1'b1;
			end
			4'b1101: begin
				correction_pattern = {4{1'b0}};correction_pattern[2]=1'b1;
			end
			4'b1110: begin
				correction_pattern = {4{1'b0}};correction_pattern[3]=1'b1;
			end
			4'b0001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b0010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b0100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b1000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_8_4_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [4-1:0] stored_data_edc = extended_hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [4-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_8_4_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_8_min_width (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_12_8_f
//Compute 4 bits Error Detection Code from a 8 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 256 valid code words out of 4096 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: x x x  x (4 inputs)
//  syndrom[1]: x  x xxx (5 inputs)
//  syndrom[2]:  xx  xxx (5 inputs)
//  syndrom[3]:  x xx x  (4 inputs)
//Input usage report:
//  input bit 0 used 2 times (syndrom bits 0 1)
//  input bit 1 used 2 times (syndrom bits 2 3)
//  input bit 2 used 2 times (syndrom bits 0 2)
//  input bit 3 used 2 times (syndrom bits 1 3)
//  input bit 4 used 2 times (syndrom bits 0 3)
//  input bit 5 used 2 times (syndrom bits 1 2)
//  input bit 6 used 3 times (syndrom bits 1 2 3)
//  input bit 7 used 3 times (syndrom bits 0 1 2)
function [4-1:0] hamming_code_12_8_f;
    input [8-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[2]^in[4]^in[7];//4 inputs
        syndrom[1] = in[0]^in[3]^in[5]^in[6]^in[7];//5 inputs
        syndrom[2] = in[1]^in[2]^in[5]^in[6]^in[7];//5 inputs
        syndrom[3] = in[1]^in[3]^in[4]^in[6];//4 inputs
        hamming_code_12_8_f = syndrom;
    end
endfunction
wire [4-1:0] stored_data_edc = hamming_code_12_8_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_8_min_width (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [5-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [5-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_13_8_f
//Compute 5 bits Error Detection Code from a 8 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 256 valid code words out of 8192 therefore 96% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: xx   xxx (5 inputs)
//  syndrom[1]: x x x xx (5 inputs)
//  syndrom[2]: x  xxx   (4 inputs)
//  syndrom[3]:  xxxx  x (5 inputs)
//  syndrom[4]:  xxx xx  (5 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 3 4)
//  input bit 2 used 3 times (syndrom bits 1 3 4)
//  input bit 3 used 3 times (syndrom bits 2 3 4)
//  input bit 4 used 3 times (syndrom bits 1 2 3)
//  input bit 5 used 3 times (syndrom bits 0 2 4)
//  input bit 6 used 3 times (syndrom bits 0 1 4)
//  input bit 7 used 3 times (syndrom bits 0 1 3)
function [5-1:0] extended_hamming_code_13_8_f;
    input [8-1:0] in;
    reg [5-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[5]^in[6]^in[7];//5 inputs
        syndrom[1] = in[0]^in[2]^in[4]^in[6]^in[7];//5 inputs
        syndrom[2] = in[0]^in[3]^in[4]^in[5];//4 inputs
        syndrom[3] = in[1]^in[2]^in[3]^in[4]^in[7];//5 inputs
        syndrom[4] = in[1]^in[2]^in[3]^in[5]^in[6];//5 inputs
        extended_hamming_code_13_8_f = syndrom;
    end
endfunction
wire [5-1:0] stored_data_edc = extended_hamming_code_13_8_f(i_stored_data);
wire [5-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_8_min_width (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [5-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [5-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [8-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_13_8_f
//Compute 5 bits Error Detection Code from a 8 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 256 valid code words out of 8192 therefore 96% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: xx   xxx (5 inputs)
//  syndrom[1]: x x x xx (5 inputs)
//  syndrom[2]: x  xxx   (4 inputs)
//  syndrom[3]:  xxxx  x (5 inputs)
//  syndrom[4]:  xxx xx  (5 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 3 4)
//  input bit 2 used 3 times (syndrom bits 1 3 4)
//  input bit 3 used 3 times (syndrom bits 2 3 4)
//  input bit 4 used 3 times (syndrom bits 1 2 3)
//  input bit 5 used 3 times (syndrom bits 0 2 4)
//  input bit 6 used 3 times (syndrom bits 0 1 4)
//  input bit 7 used 3 times (syndrom bits 0 1 3)
function [5-1:0] extended_hamming_code_13_8_f;
    input [8-1:0] in;
    reg [5-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[5]^in[6]^in[7];//5 inputs
        syndrom[1] = in[0]^in[2]^in[4]^in[6]^in[7];//5 inputs
        syndrom[2] = in[0]^in[3]^in[4]^in[5];//4 inputs
        syndrom[3] = in[1]^in[2]^in[3]^in[4]^in[7];//5 inputs
        syndrom[4] = in[1]^in[2]^in[3]^in[5]^in[6];//5 inputs
        extended_hamming_code_13_8_f = syndrom;
    end
endfunction
function [2+8-1:0] extended_hamming_code_13_8_f_correction_pattern_f;
    input [5-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [8-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {8{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			5'b00000: begin
				correctable_error = 1'b0;
				correction_pattern = {8{1'b0}};
			end	
			5'b00111: begin
				correction_pattern = {8{1'b0}};correction_pattern[0]=1'b1;
			end
			5'b11001: begin
				correction_pattern = {8{1'b0}};correction_pattern[1]=1'b1;
			end
			5'b11010: begin
				correction_pattern = {8{1'b0}};correction_pattern[2]=1'b1;
			end
			5'b11100: begin
				correction_pattern = {8{1'b0}};correction_pattern[3]=1'b1;
			end
			5'b01110: begin
				correction_pattern = {8{1'b0}};correction_pattern[4]=1'b1;
			end
			5'b10101: begin
				correction_pattern = {8{1'b0}};correction_pattern[5]=1'b1;
			end
			5'b10011: begin
				correction_pattern = {8{1'b0}};correction_pattern[6]=1'b1;
			end
			5'b01011: begin
				correction_pattern = {8{1'b0}};correction_pattern[7]=1'b1;
			end
			5'b00001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			5'b00010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			5'b00100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			5'b01000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			5'b10000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_13_8_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [5-1:0] stored_data_edc = extended_hamming_code_13_8_f(i_stored_data);
wire [5-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [8-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_13_8_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_12_min_width (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [5-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [5-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_17_12_f
//Compute 5 bits Error Detection Code from a 12 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 131072 therefore 96% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[0]: x   x  xx x  (5 inputs)
//  syndrom[1]: x    xx  xxx (6 inputs)
//  syndrom[2]:  xx   xx   x (5 inputs)
//  syndrom[3]:  x x x  x  x (5 inputs)
//  syndrom[4]:   xxx    xx  (5 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 2 4)
//  input bit  3 used 2 times (syndrom bits 3 4)
//  input bit  4 used 2 times (syndrom bits 0 4)
//  input bit  5 used 2 times (syndrom bits 1 3)
//  input bit  6 used 2 times (syndrom bits 1 2)
//  input bit  7 used 2 times (syndrom bits 0 2)
//  input bit  8 used 2 times (syndrom bits 0 3)
//  input bit  9 used 2 times (syndrom bits 1 4)
//  input bit 10 used 3 times (syndrom bits 0 1 4)
//  input bit 11 used 3 times (syndrom bits 1 2 3)
function [5-1:0] hamming_code_17_12_f;
    input [12-1:0] in;
    reg [5-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 7]^in[ 8]^in[10];//5 inputs
        syndrom[1] = in[ 0]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[11];//6 inputs
        syndrom[2] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[11];//5 inputs
        syndrom[3] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[11];//5 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10];//5 inputs
        hamming_code_17_12_f = syndrom;
    end
endfunction
wire [5-1:0] stored_data_edc = hamming_code_17_12_f(i_stored_data);
wire [5-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_12_min_width (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_18_12_f
//Compute 6 bits Error Detection Code from a 12 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 262144 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[0]: x x  x xx x  (6 inputs)
//  syndrom[1]: x  xx  xx  x (6 inputs)
//  syndrom[2]: x  x xx  xx  (6 inputs)
//  syndrom[3]:  xx x  x xx  (6 inputs)
//  syndrom[4]:  xx  xx x  x (6 inputs)
//  syndrom[5]:  x xx x  x x (6 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
function [6-1:0] extended_hamming_code_18_12_f;
    input [12-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10];//6 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11];//6 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10];//6 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10];//6 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11];//6 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11];//6 inputs
        extended_hamming_code_18_12_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = extended_hamming_code_18_12_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_12_min_width (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [12-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_18_12_f
//Compute 6 bits Error Detection Code from a 12 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 262144 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[0]: x x  x xx x  (6 inputs)
//  syndrom[1]: x  xx  xx  x (6 inputs)
//  syndrom[2]: x  x xx  xx  (6 inputs)
//  syndrom[3]:  xx x  x xx  (6 inputs)
//  syndrom[4]:  xx  xx x  x (6 inputs)
//  syndrom[5]:  x xx x  x x (6 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
function [6-1:0] extended_hamming_code_18_12_f;
    input [12-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10];//6 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11];//6 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10];//6 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10];//6 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11];//6 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11];//6 inputs
        extended_hamming_code_18_12_f = syndrom;
    end
endfunction
function [2+12-1:0] extended_hamming_code_18_12_f_correction_pattern_f;
    input [6-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [12-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {12{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			6'b000000: begin
				correctable_error = 1'b0;
				correction_pattern = {12{1'b0}};
			end	
			6'b000111: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 0]=1'b1;
			end
			6'b111000: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 1]=1'b1;
			end
			6'b011001: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 2]=1'b1;
			end
			6'b100110: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 3]=1'b1;
			end
			6'b101010: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 4]=1'b1;
			end
			6'b010101: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 5]=1'b1;
			end
			6'b110100: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 6]=1'b1;
			end
			6'b001011: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 7]=1'b1;
			end
			6'b010011: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 8]=1'b1;
			end
			6'b101100: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 9]=1'b1;
			end
			6'b001101: begin
				correction_pattern = {12{1'b0}};correction_pattern[10]=1'b1;
			end
			6'b110010: begin
				correction_pattern = {12{1'b0}};correction_pattern[11]=1'b1;
			end
			6'b000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_18_12_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [6-1:0] stored_data_edc = extended_hamming_code_18_12_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [12-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_18_12_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_16_min_width (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [5-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [5-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_21_16_f
//Compute 5 bits Error Detection Code from a 16 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 2097152 therefore 96% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[0]: x   x  xx x  xxx (8 inputs)
//  syndrom[1]: x    xx  xxx   x (7 inputs)
//  syndrom[2]:  xx   xx   xxx x (8 inputs)
//  syndrom[3]:  x x x  x  xxxx  (8 inputs)
//  syndrom[4]:   xxx    xx x x  (7 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 2 4)
//  input bit  3 used 2 times (syndrom bits 3 4)
//  input bit  4 used 2 times (syndrom bits 0 4)
//  input bit  5 used 2 times (syndrom bits 1 3)
//  input bit  6 used 2 times (syndrom bits 1 2)
//  input bit  7 used 2 times (syndrom bits 0 2)
//  input bit  8 used 2 times (syndrom bits 0 3)
//  input bit  9 used 2 times (syndrom bits 1 4)
//  input bit 10 used 3 times (syndrom bits 0 1 4)
//  input bit 11 used 3 times (syndrom bits 1 2 3)
//  input bit 12 used 3 times (syndrom bits 2 3 4)
//  input bit 13 used 3 times (syndrom bits 0 2 3)
//  input bit 14 used 3 times (syndrom bits 0 3 4)
//  input bit 15 used 3 times (syndrom bits 0 1 2)
function [5-1:0] hamming_code_21_16_f;
    input [16-1:0] in;
    reg [5-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 7]^in[ 8]^in[10]^in[13]^in[14]^in[15];//8 inputs
        syndrom[1] = in[ 0]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[11]^in[15];//7 inputs
        syndrom[2] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[11]^in[12]^in[13]^in[15];//8 inputs
        syndrom[3] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[11]^in[12]^in[13]^in[14];//8 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[12]^in[14];//7 inputs
        hamming_code_21_16_f = syndrom;
    end
endfunction
wire [5-1:0] stored_data_edc = hamming_code_21_16_f(i_stored_data);
wire [5-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_16_min_width (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_22_16_f
//Compute 6 bits Error Detection Code from a 16 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 4194304 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[0]: x x  x xx x x  x (8 inputs)
//  syndrom[1]: x  xx  xx  xx x  (8 inputs)
//  syndrom[2]: x  x xx  xx  x x (8 inputs)
//  syndrom[3]:  xx x  x xx  xx  (8 inputs)
//  syndrom[4]:  xx  xx x  x xx  (8 inputs)
//  syndrom[5]:  x xx x  x xx  x (8 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
function [6-1:0] extended_hamming_code_22_16_f;
    input [16-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10]^in[12]^in[15];//8 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11]^in[12]^in[14];//8 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[13]^in[15];//8 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10]^in[13]^in[14];//8 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11]^in[13]^in[14];//8 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11]^in[12]^in[15];//8 inputs
        extended_hamming_code_22_16_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = extended_hamming_code_22_16_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_16_min_width (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [16-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_22_16_f
//Compute 6 bits Error Detection Code from a 16 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 4194304 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[0]: x x  x xx x x  x (8 inputs)
//  syndrom[1]: x  xx  xx  xx x  (8 inputs)
//  syndrom[2]: x  x xx  xx  x x (8 inputs)
//  syndrom[3]:  xx x  x xx  xx  (8 inputs)
//  syndrom[4]:  xx  xx x  x xx  (8 inputs)
//  syndrom[5]:  x xx x  x xx  x (8 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
function [6-1:0] extended_hamming_code_22_16_f;
    input [16-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10]^in[12]^in[15];//8 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11]^in[12]^in[14];//8 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[13]^in[15];//8 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10]^in[13]^in[14];//8 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11]^in[13]^in[14];//8 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11]^in[12]^in[15];//8 inputs
        extended_hamming_code_22_16_f = syndrom;
    end
endfunction
function [2+16-1:0] extended_hamming_code_22_16_f_correction_pattern_f;
    input [6-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [16-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {16{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			6'b000000: begin
				correctable_error = 1'b0;
				correction_pattern = {16{1'b0}};
			end	
			6'b000111: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 0]=1'b1;
			end
			6'b111000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 1]=1'b1;
			end
			6'b011001: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 2]=1'b1;
			end
			6'b100110: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 3]=1'b1;
			end
			6'b101010: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 4]=1'b1;
			end
			6'b010101: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 5]=1'b1;
			end
			6'b110100: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 6]=1'b1;
			end
			6'b001011: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 7]=1'b1;
			end
			6'b010011: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 8]=1'b1;
			end
			6'b101100: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 9]=1'b1;
			end
			6'b001101: begin
				correction_pattern = {16{1'b0}};correction_pattern[10]=1'b1;
			end
			6'b110010: begin
				correction_pattern = {16{1'b0}};correction_pattern[11]=1'b1;
			end
			6'b100011: begin
				correction_pattern = {16{1'b0}};correction_pattern[12]=1'b1;
			end
			6'b011100: begin
				correction_pattern = {16{1'b0}};correction_pattern[13]=1'b1;
			end
			6'b011010: begin
				correction_pattern = {16{1'b0}};correction_pattern[14]=1'b1;
			end
			6'b100101: begin
				correction_pattern = {16{1'b0}};correction_pattern[15]=1'b1;
			end
			6'b000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_22_16_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [6-1:0] stored_data_edc = extended_hamming_code_22_16_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [16-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_22_16_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_20_min_width (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [5-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [5-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_25_20_f
//Compute 5 bits Error Detection Code from a 20 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 33554432 therefore 96% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[0]: x   x  xx x  xxx  xx (10 inputs)
//  syndrom[1]: x    xx  xxx   xxxx  (10 inputs)
//  syndrom[2]:  xx   xx   xxx xx  x (10 inputs)
//  syndrom[3]:  x x x  x  xxxx  xx  (10 inputs)
//  syndrom[4]:   xxx    xx x x xx x (10 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 2 4)
//  input bit  3 used 2 times (syndrom bits 3 4)
//  input bit  4 used 2 times (syndrom bits 0 4)
//  input bit  5 used 2 times (syndrom bits 1 3)
//  input bit  6 used 2 times (syndrom bits 1 2)
//  input bit  7 used 2 times (syndrom bits 0 2)
//  input bit  8 used 2 times (syndrom bits 0 3)
//  input bit  9 used 2 times (syndrom bits 1 4)
//  input bit 10 used 3 times (syndrom bits 0 1 4)
//  input bit 11 used 3 times (syndrom bits 1 2 3)
//  input bit 12 used 3 times (syndrom bits 2 3 4)
//  input bit 13 used 3 times (syndrom bits 0 2 3)
//  input bit 14 used 3 times (syndrom bits 0 3 4)
//  input bit 15 used 3 times (syndrom bits 0 1 2)
//  input bit 16 used 3 times (syndrom bits 1 2 4)
//  input bit 17 used 3 times (syndrom bits 1 3 4)
//  input bit 18 used 3 times (syndrom bits 0 1 3)
//  input bit 19 used 3 times (syndrom bits 0 2 4)
function [5-1:0] hamming_code_25_20_f;
    input [20-1:0] in;
    reg [5-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 7]^in[ 8]^in[10]^in[13]^in[14]^in[15]^in[18]^in[19];//10 inputs
        syndrom[1] = in[ 0]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[11]^in[15]^in[16]^in[17]^in[18];//10 inputs
        syndrom[2] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[11]^in[12]^in[13]^in[15]^in[16]^in[19];//10 inputs
        syndrom[3] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[11]^in[12]^in[13]^in[14]^in[17]^in[18];//10 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[12]^in[14]^in[16]^in[17]^in[19];//10 inputs
        hamming_code_25_20_f = syndrom;
    end
endfunction
wire [5-1:0] stored_data_edc = hamming_code_25_20_f(i_stored_data);
wire [5-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_20_min_width (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_26_20_f
//Compute 6 bits Error Detection Code from a 20 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 67108864 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[0]: x x  x xx x x  x xx  (10 inputs)
//  syndrom[1]: x  xx  xx  xx x x  x (10 inputs)
//  syndrom[2]: x  x xx  xx  x xx  x (10 inputs)
//  syndrom[3]:  xx x  x xx  xx  x x (10 inputs)
//  syndrom[4]:  xx  xx x  x xx x x  (10 inputs)
//  syndrom[5]:  x xx x  x xx  x xx  (10 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 1 2 4)
//  input bit 17 used 3 times (syndrom bits 0 3 5)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 1 2 3)
function [6-1:0] extended_hamming_code_26_20_f;
    input [20-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[18];//10 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11]^in[12]^in[14]^in[16]^in[19];//10 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[13]^in[15]^in[16]^in[19];//10 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10]^in[13]^in[14]^in[17]^in[19];//10 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11]^in[13]^in[14]^in[16]^in[18];//10 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11]^in[12]^in[15]^in[17]^in[18];//10 inputs
        extended_hamming_code_26_20_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = extended_hamming_code_26_20_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_20_min_width (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [20-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_26_20_f
//Compute 6 bits Error Detection Code from a 20 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 67108864 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[0]: x x  x xx x x  x xx  (10 inputs)
//  syndrom[1]: x  xx  xx  xx x x  x (10 inputs)
//  syndrom[2]: x  x xx  xx  x xx  x (10 inputs)
//  syndrom[3]:  xx x  x xx  xx  x x (10 inputs)
//  syndrom[4]:  xx  xx x  x xx x x  (10 inputs)
//  syndrom[5]:  x xx x  x xx  x xx  (10 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 1 2 4)
//  input bit 17 used 3 times (syndrom bits 0 3 5)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 1 2 3)
function [6-1:0] extended_hamming_code_26_20_f;
    input [20-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[18];//10 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11]^in[12]^in[14]^in[16]^in[19];//10 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[13]^in[15]^in[16]^in[19];//10 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10]^in[13]^in[14]^in[17]^in[19];//10 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11]^in[13]^in[14]^in[16]^in[18];//10 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11]^in[12]^in[15]^in[17]^in[18];//10 inputs
        extended_hamming_code_26_20_f = syndrom;
    end
endfunction
function [2+20-1:0] extended_hamming_code_26_20_f_correction_pattern_f;
    input [6-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [20-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {20{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			6'b000000: begin
				correctable_error = 1'b0;
				correction_pattern = {20{1'b0}};
			end	
			6'b000111: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 0]=1'b1;
			end
			6'b111000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 1]=1'b1;
			end
			6'b011001: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 2]=1'b1;
			end
			6'b100110: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 3]=1'b1;
			end
			6'b101010: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 4]=1'b1;
			end
			6'b010101: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 5]=1'b1;
			end
			6'b110100: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 6]=1'b1;
			end
			6'b001011: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 7]=1'b1;
			end
			6'b010011: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 8]=1'b1;
			end
			6'b101100: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 9]=1'b1;
			end
			6'b001101: begin
				correction_pattern = {20{1'b0}};correction_pattern[10]=1'b1;
			end
			6'b110010: begin
				correction_pattern = {20{1'b0}};correction_pattern[11]=1'b1;
			end
			6'b100011: begin
				correction_pattern = {20{1'b0}};correction_pattern[12]=1'b1;
			end
			6'b011100: begin
				correction_pattern = {20{1'b0}};correction_pattern[13]=1'b1;
			end
			6'b011010: begin
				correction_pattern = {20{1'b0}};correction_pattern[14]=1'b1;
			end
			6'b100101: begin
				correction_pattern = {20{1'b0}};correction_pattern[15]=1'b1;
			end
			6'b010110: begin
				correction_pattern = {20{1'b0}};correction_pattern[16]=1'b1;
			end
			6'b101001: begin
				correction_pattern = {20{1'b0}};correction_pattern[17]=1'b1;
			end
			6'b110001: begin
				correction_pattern = {20{1'b0}};correction_pattern[18]=1'b1;
			end
			6'b001110: begin
				correction_pattern = {20{1'b0}};correction_pattern[19]=1'b1;
			end
			6'b000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_26_20_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [6-1:0] stored_data_edc = extended_hamming_code_26_20_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [20-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_26_20_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_24_min_width (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [5-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [5-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_29_24_f
//Compute 5 bits Error Detection Code from a 24 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 536870912 therefore 96% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[0]: x   x  xx x  xxx  xxxxxx (14 inputs)
//  syndrom[1]: x    xx  xxx   xxxx x xx (13 inputs)
//  syndrom[2]:  xx   xx   xxx xx  xxx x (13 inputs)
//  syndrom[3]:  x x x  x  xxxx  xx  xxx (13 inputs)
//  syndrom[4]:   xxx    xx x x xx xxxx  (13 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 2 4)
//  input bit  3 used 2 times (syndrom bits 3 4)
//  input bit  4 used 2 times (syndrom bits 0 4)
//  input bit  5 used 2 times (syndrom bits 1 3)
//  input bit  6 used 2 times (syndrom bits 1 2)
//  input bit  7 used 2 times (syndrom bits 0 2)
//  input bit  8 used 2 times (syndrom bits 0 3)
//  input bit  9 used 2 times (syndrom bits 1 4)
//  input bit 10 used 3 times (syndrom bits 0 1 4)
//  input bit 11 used 3 times (syndrom bits 1 2 3)
//  input bit 12 used 3 times (syndrom bits 2 3 4)
//  input bit 13 used 3 times (syndrom bits 0 2 3)
//  input bit 14 used 3 times (syndrom bits 0 3 4)
//  input bit 15 used 3 times (syndrom bits 0 1 2)
//  input bit 16 used 3 times (syndrom bits 1 2 4)
//  input bit 17 used 3 times (syndrom bits 1 3 4)
//  input bit 18 used 3 times (syndrom bits 0 1 3)
//  input bit 19 used 3 times (syndrom bits 0 2 4)
//  input bit 20 used 4 times (syndrom bits 0 1 2 4)
//  input bit 21 used 4 times (syndrom bits 0 2 3 4)
//  input bit 22 used 4 times (syndrom bits 0 1 3 4)
//  input bit 23 used 4 times (syndrom bits 0 1 2 3)
function [5-1:0] hamming_code_29_24_f;
    input [24-1:0] in;
    reg [5-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 7]^in[ 8]^in[10]^in[13]^in[14]^in[15]^in[18]^in[19]^in[20]^in[21]^in[22]^in[23];//14 inputs
        syndrom[1] = in[ 0]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[11]^in[15]^in[16]^in[17]^in[18]^in[20]^in[22]^in[23];//13 inputs
        syndrom[2] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[11]^in[12]^in[13]^in[15]^in[16]^in[19]^in[20]^in[21]^in[23];//13 inputs
        syndrom[3] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[11]^in[12]^in[13]^in[14]^in[17]^in[18]^in[21]^in[22]^in[23];//13 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[12]^in[14]^in[16]^in[17]^in[19]^in[20]^in[21]^in[22];//13 inputs
        hamming_code_29_24_f = syndrom;
    end
endfunction
wire [5-1:0] stored_data_edc = hamming_code_29_24_f(i_stored_data);
wire [5-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_24_min_width (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_30_24_f
//Compute 6 bits Error Detection Code from a 24 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 1073741824 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[0]: x x  x xx x x  x xx x xx (13 inputs)
//  syndrom[1]: x  xx  xx  xx x x  xxxx  (13 inputs)
//  syndrom[2]: x  x xx  xx  x xx  xxxxx (14 inputs)
//  syndrom[3]:  xx x  x xx  xx  x xxxxx (14 inputs)
//  syndrom[4]:  xx  xx x  x xx x x  xxx (13 inputs)
//  syndrom[5]:  x xx x  x xx  x xx xx x (13 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 1 2 4)
//  input bit 17 used 3 times (syndrom bits 0 3 5)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 1 2 3)
//  input bit 20 used 5 times (syndrom bits 0 1 2 3 5)
//  input bit 21 used 5 times (syndrom bits 1 2 3 4 5)
//  input bit 22 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 23 used 5 times (syndrom bits 0 2 3 4 5)
function [6-1:0] extended_hamming_code_30_24_f;
    input [24-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[18]^in[20]^in[22]^in[23];//13 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11]^in[12]^in[14]^in[16]^in[19]^in[20]^in[21]^in[22];//13 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[13]^in[15]^in[16]^in[19]^in[20]^in[21]^in[22]^in[23];//14 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10]^in[13]^in[14]^in[17]^in[19]^in[20]^in[21]^in[22]^in[23];//14 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11]^in[13]^in[14]^in[16]^in[18]^in[21]^in[22]^in[23];//13 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11]^in[12]^in[15]^in[17]^in[18]^in[20]^in[21]^in[23];//13 inputs
        extended_hamming_code_30_24_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = extended_hamming_code_30_24_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_24_min_width (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [24-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_30_24_f
//Compute 6 bits Error Detection Code from a 24 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 1073741824 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[0]: x x  x xx x x  x xx x xx (13 inputs)
//  syndrom[1]: x  xx  xx  xx x x  xxxx  (13 inputs)
//  syndrom[2]: x  x xx  xx  x xx  xxxxx (14 inputs)
//  syndrom[3]:  xx x  x xx  xx  x xxxxx (14 inputs)
//  syndrom[4]:  xx  xx x  x xx x x  xxx (13 inputs)
//  syndrom[5]:  x xx x  x xx  x xx xx x (13 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 1 2 4)
//  input bit 17 used 3 times (syndrom bits 0 3 5)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 1 2 3)
//  input bit 20 used 5 times (syndrom bits 0 1 2 3 5)
//  input bit 21 used 5 times (syndrom bits 1 2 3 4 5)
//  input bit 22 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 23 used 5 times (syndrom bits 0 2 3 4 5)
function [6-1:0] extended_hamming_code_30_24_f;
    input [24-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[18]^in[20]^in[22]^in[23];//13 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11]^in[12]^in[14]^in[16]^in[19]^in[20]^in[21]^in[22];//13 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10]^in[13]^in[15]^in[16]^in[19]^in[20]^in[21]^in[22]^in[23];//14 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10]^in[13]^in[14]^in[17]^in[19]^in[20]^in[21]^in[22]^in[23];//14 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11]^in[13]^in[14]^in[16]^in[18]^in[21]^in[22]^in[23];//13 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11]^in[12]^in[15]^in[17]^in[18]^in[20]^in[21]^in[23];//13 inputs
        extended_hamming_code_30_24_f = syndrom;
    end
endfunction
function [2+24-1:0] extended_hamming_code_30_24_f_correction_pattern_f;
    input [6-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [24-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {24{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			6'b000000: begin
				correctable_error = 1'b0;
				correction_pattern = {24{1'b0}};
			end	
			6'b000111: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 0]=1'b1;
			end
			6'b111000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 1]=1'b1;
			end
			6'b011001: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 2]=1'b1;
			end
			6'b100110: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 3]=1'b1;
			end
			6'b101010: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 4]=1'b1;
			end
			6'b010101: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 5]=1'b1;
			end
			6'b110100: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 6]=1'b1;
			end
			6'b001011: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 7]=1'b1;
			end
			6'b010011: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 8]=1'b1;
			end
			6'b101100: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 9]=1'b1;
			end
			6'b001101: begin
				correction_pattern = {24{1'b0}};correction_pattern[10]=1'b1;
			end
			6'b110010: begin
				correction_pattern = {24{1'b0}};correction_pattern[11]=1'b1;
			end
			6'b100011: begin
				correction_pattern = {24{1'b0}};correction_pattern[12]=1'b1;
			end
			6'b011100: begin
				correction_pattern = {24{1'b0}};correction_pattern[13]=1'b1;
			end
			6'b011010: begin
				correction_pattern = {24{1'b0}};correction_pattern[14]=1'b1;
			end
			6'b100101: begin
				correction_pattern = {24{1'b0}};correction_pattern[15]=1'b1;
			end
			6'b010110: begin
				correction_pattern = {24{1'b0}};correction_pattern[16]=1'b1;
			end
			6'b101001: begin
				correction_pattern = {24{1'b0}};correction_pattern[17]=1'b1;
			end
			6'b110001: begin
				correction_pattern = {24{1'b0}};correction_pattern[18]=1'b1;
			end
			6'b001110: begin
				correction_pattern = {24{1'b0}};correction_pattern[19]=1'b1;
			end
			6'b101111: begin
				correction_pattern = {24{1'b0}};correction_pattern[20]=1'b1;
			end
			6'b111110: begin
				correction_pattern = {24{1'b0}};correction_pattern[21]=1'b1;
			end
			6'b011111: begin
				correction_pattern = {24{1'b0}};correction_pattern[22]=1'b1;
			end
			6'b111101: begin
				correction_pattern = {24{1'b0}};correction_pattern[23]=1'b1;
			end
			6'b000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_30_24_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [6-1:0] stored_data_edc = extended_hamming_code_30_24_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [24-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_30_24_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_32_min_width (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_38_32_f
//Compute 6 bits Error Detection Code from a 32 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 274877906944 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[0]: x    x  xx x    x xx x  x xx  x  (13 inputs)
//  syndrom[1]: x     xx  x  x  xx x  x xx  xx   (13 inputs)
//  syndrom[2]:  x x    x x x   xx  xx x  x xx x (14 inputs)
//  syndrom[3]:  x  x x    x  xx x  x xx x x  x  (13 inputs)
//  syndrom[4]:   xx   x x    xx  xx  xx  xx x x (14 inputs)
//  syndrom[5]:   x xx      xx x  x xx  xx  x xx (14 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 2 4)
//  input bit  4 used 2 times (syndrom bits 3 5)
//  input bit  5 used 2 times (syndrom bits 0 5)
//  input bit  6 used 2 times (syndrom bits 1 3)
//  input bit  7 used 2 times (syndrom bits 1 4)
//  input bit  8 used 2 times (syndrom bits 0 2)
//  input bit  9 used 2 times (syndrom bits 0 4)
//  input bit 10 used 2 times (syndrom bits 1 2)
//  input bit 11 used 2 times (syndrom bits 0 3)
//  input bit 12 used 2 times (syndrom bits 2 5)
//  input bit 13 used 2 times (syndrom bits 1 5)
//  input bit 14 used 2 times (syndrom bits 3 4)
//  input bit 15 used 3 times (syndrom bits 3 4 5)
//  input bit 16 used 3 times (syndrom bits 0 1 2)
//  input bit 17 used 3 times (syndrom bits 1 2 3)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 0 1 4)
//  input bit 20 used 3 times (syndrom bits 2 3 5)
//  input bit 21 used 3 times (syndrom bits 0 2 5)
//  input bit 22 used 3 times (syndrom bits 1 3 4)
//  input bit 23 used 3 times (syndrom bits 2 3 4)
//  input bit 24 used 3 times (syndrom bits 0 1 5)
//  input bit 25 used 3 times (syndrom bits 1 3 5)
//  input bit 26 used 3 times (syndrom bits 0 2 4)
//  input bit 27 used 3 times (syndrom bits 0 3 4)
//  input bit 28 used 3 times (syndrom bits 1 2 5)
//  input bit 29 used 3 times (syndrom bits 1 2 4)
//  input bit 30 used 3 times (syndrom bits 0 3 5)
//  input bit 31 used 3 times (syndrom bits 2 4 5)
function [6-1:0] hamming_code_38_32_f;
    input [32-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 5]^in[ 8]^in[ 9]^in[11]^in[16]^in[18]^in[19]^in[21]^in[24]^in[26]^in[27]^in[30];//13 inputs
        syndrom[1] = in[ 0]^in[ 6]^in[ 7]^in[10]^in[13]^in[16]^in[17]^in[19]^in[22]^in[24]^in[25]^in[28]^in[29];//13 inputs
        syndrom[2] = in[ 1]^in[ 3]^in[ 8]^in[10]^in[12]^in[16]^in[17]^in[20]^in[21]^in[23]^in[26]^in[28]^in[29]^in[31];//14 inputs
        syndrom[3] = in[ 1]^in[ 4]^in[ 6]^in[11]^in[14]^in[15]^in[17]^in[20]^in[22]^in[23]^in[25]^in[27]^in[30];//13 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 7]^in[ 9]^in[14]^in[15]^in[18]^in[19]^in[22]^in[23]^in[26]^in[27]^in[29]^in[31];//14 inputs
        syndrom[5] = in[ 2]^in[ 4]^in[ 5]^in[12]^in[13]^in[15]^in[18]^in[20]^in[21]^in[24]^in[25]^in[28]^in[30]^in[31];//14 inputs
        hamming_code_38_32_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = hamming_code_38_32_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_32_min_width (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_39_32_f
//Compute 7 bits Error Detection Code from a 32 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 549755813888 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx  (14 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x (14 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx    (13 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx    (13 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx  (14 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x (14 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xx (14 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
function [7-1:0] extended_hamming_code_39_32_f;
    input [32-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30];//14 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31];//14 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28];//13 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28];//13 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30];//14 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31];//14 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31];//14 inputs
        extended_hamming_code_39_32_f = syndrom;
    end
endfunction
wire [7-1:0] stored_data_edc = extended_hamming_code_39_32_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_32_min_width (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [32-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_39_32_f
//Compute 7 bits Error Detection Code from a 32 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 549755813888 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx  (14 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x (14 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx    (13 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx    (13 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx  (14 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x (14 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xx (14 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
function [7-1:0] extended_hamming_code_39_32_f;
    input [32-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30];//14 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31];//14 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28];//13 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28];//13 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30];//14 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31];//14 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31];//14 inputs
        extended_hamming_code_39_32_f = syndrom;
    end
endfunction
function [2+32-1:0] extended_hamming_code_39_32_f_correction_pattern_f;
    input [7-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [32-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {32{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			7'b0000000: begin
				correctable_error = 1'b0;
				correction_pattern = {32{1'b0}};
			end	
			7'b0000111: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 0]=1'b1;
			end
			7'b0111000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 1]=1'b1;
			end
			7'b1011000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 2]=1'b1;
			end
			7'b1100001: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 3]=1'b1;
			end
			7'b1000110: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 4]=1'b1;
			end
			7'b0100110: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 5]=1'b1;
			end
			7'b0011001: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 6]=1'b1;
			end
			7'b0001011: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 7]=1'b1;
			end
			7'b0110100: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 8]=1'b1;
			end
			7'b1010100: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 9]=1'b1;
			end
			7'b1101000: begin
				correction_pattern = {32{1'b0}};correction_pattern[10]=1'b1;
			end
			7'b1000011: begin
				correction_pattern = {32{1'b0}};correction_pattern[11]=1'b1;
			end
			7'b0100011: begin
				correction_pattern = {32{1'b0}};correction_pattern[12]=1'b1;
			end
			7'b0011100: begin
				correction_pattern = {32{1'b0}};correction_pattern[13]=1'b1;
			end
			7'b0011010: begin
				correction_pattern = {32{1'b0}};correction_pattern[14]=1'b1;
			end
			7'b0100101: begin
				correction_pattern = {32{1'b0}};correction_pattern[15]=1'b1;
			end
			7'b1000101: begin
				correction_pattern = {32{1'b0}};correction_pattern[16]=1'b1;
			end
			7'b1110000: begin
				correction_pattern = {32{1'b0}};correction_pattern[17]=1'b1;
			end
			7'b1001010: begin
				correction_pattern = {32{1'b0}};correction_pattern[18]=1'b1;
			end
			7'b0101010: begin
				correction_pattern = {32{1'b0}};correction_pattern[19]=1'b1;
			end
			7'b0010101: begin
				correction_pattern = {32{1'b0}};correction_pattern[20]=1'b1;
			end
			7'b0010110: begin
				correction_pattern = {32{1'b0}};correction_pattern[21]=1'b1;
			end
			7'b0101001: begin
				correction_pattern = {32{1'b0}};correction_pattern[22]=1'b1;
			end
			7'b1001001: begin
				correction_pattern = {32{1'b0}};correction_pattern[23]=1'b1;
			end
			7'b1100100: begin
				correction_pattern = {32{1'b0}};correction_pattern[24]=1'b1;
			end
			7'b1010010: begin
				correction_pattern = {32{1'b0}};correction_pattern[25]=1'b1;
			end
			7'b0110010: begin
				correction_pattern = {32{1'b0}};correction_pattern[26]=1'b1;
			end
			7'b0001101: begin
				correction_pattern = {32{1'b0}};correction_pattern[27]=1'b1;
			end
			7'b0001110: begin
				correction_pattern = {32{1'b0}};correction_pattern[28]=1'b1;
			end
			7'b0110001: begin
				correction_pattern = {32{1'b0}};correction_pattern[29]=1'b1;
			end
			7'b1010001: begin
				correction_pattern = {32{1'b0}};correction_pattern[30]=1'b1;
			end
			7'b1100010: begin
				correction_pattern = {32{1'b0}};correction_pattern[31]=1'b1;
			end
			7'b0000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b1000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_39_32_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [7-1:0] stored_data_edc = extended_hamming_code_39_32_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [32-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_39_32_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_36_min_width (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_42_36_f
//Compute 6 bits Error Detection Code from a 36 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 4398046511104 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[0]: x    x  xx x    x xx x  x xx  x xx x (16 inputs)
//  syndrom[1]: x     xx  x  x  xx x  x xx  xx  x xx (16 inputs)
//  syndrom[2]:  x x    x x x   xx  xx x  x xx x x   (15 inputs)
//  syndrom[3]:  x  x x    x  xx x  x xx x x  x xx   (15 inputs)
//  syndrom[4]:   xx   x x    xx  xx  xx  xx x x  xx (16 inputs)
//  syndrom[5]:   x xx      xx x  x xx  xx  x xx  xx (16 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 2 4)
//  input bit  4 used 2 times (syndrom bits 3 5)
//  input bit  5 used 2 times (syndrom bits 0 5)
//  input bit  6 used 2 times (syndrom bits 1 3)
//  input bit  7 used 2 times (syndrom bits 1 4)
//  input bit  8 used 2 times (syndrom bits 0 2)
//  input bit  9 used 2 times (syndrom bits 0 4)
//  input bit 10 used 2 times (syndrom bits 1 2)
//  input bit 11 used 2 times (syndrom bits 0 3)
//  input bit 12 used 2 times (syndrom bits 2 5)
//  input bit 13 used 2 times (syndrom bits 1 5)
//  input bit 14 used 2 times (syndrom bits 3 4)
//  input bit 15 used 3 times (syndrom bits 3 4 5)
//  input bit 16 used 3 times (syndrom bits 0 1 2)
//  input bit 17 used 3 times (syndrom bits 1 2 3)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 0 1 4)
//  input bit 20 used 3 times (syndrom bits 2 3 5)
//  input bit 21 used 3 times (syndrom bits 0 2 5)
//  input bit 22 used 3 times (syndrom bits 1 3 4)
//  input bit 23 used 3 times (syndrom bits 2 3 4)
//  input bit 24 used 3 times (syndrom bits 0 1 5)
//  input bit 25 used 3 times (syndrom bits 1 3 5)
//  input bit 26 used 3 times (syndrom bits 0 2 4)
//  input bit 27 used 3 times (syndrom bits 0 3 4)
//  input bit 28 used 3 times (syndrom bits 1 2 5)
//  input bit 29 used 3 times (syndrom bits 1 2 4)
//  input bit 30 used 3 times (syndrom bits 0 3 5)
//  input bit 31 used 3 times (syndrom bits 2 4 5)
//  input bit 32 used 3 times (syndrom bits 0 1 3)
//  input bit 33 used 3 times (syndrom bits 0 2 3)
//  input bit 34 used 3 times (syndrom bits 1 4 5)
//  input bit 35 used 4 times (syndrom bits 0 1 4 5)
function [6-1:0] hamming_code_42_36_f;
    input [36-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 5]^in[ 8]^in[ 9]^in[11]^in[16]^in[18]^in[19]^in[21]^in[24]^in[26]^in[27]^in[30]^in[32]^in[33]^in[35];//16 inputs
        syndrom[1] = in[ 0]^in[ 6]^in[ 7]^in[10]^in[13]^in[16]^in[17]^in[19]^in[22]^in[24]^in[25]^in[28]^in[29]^in[32]^in[34]^in[35];//16 inputs
        syndrom[2] = in[ 1]^in[ 3]^in[ 8]^in[10]^in[12]^in[16]^in[17]^in[20]^in[21]^in[23]^in[26]^in[28]^in[29]^in[31]^in[33];//15 inputs
        syndrom[3] = in[ 1]^in[ 4]^in[ 6]^in[11]^in[14]^in[15]^in[17]^in[20]^in[22]^in[23]^in[25]^in[27]^in[30]^in[32]^in[33];//15 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 7]^in[ 9]^in[14]^in[15]^in[18]^in[19]^in[22]^in[23]^in[26]^in[27]^in[29]^in[31]^in[34]^in[35];//16 inputs
        syndrom[5] = in[ 2]^in[ 4]^in[ 5]^in[12]^in[13]^in[15]^in[18]^in[20]^in[21]^in[24]^in[25]^in[28]^in[30]^in[31]^in[34]^in[35];//16 inputs
        hamming_code_42_36_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = hamming_code_42_36_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_36_min_width (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_43_36_f
//Compute 7 bits Error Detection Code from a 36 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 8796093022208 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx   xx (16 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x  xx (16 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx   xx x (16 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx   xx x (16 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx   xx (16 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x x   (15 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xxx    (15 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
//  input bit 32 used 3 times (syndrom bits 2 3 6)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 1 4)
//  input bit 35 used 5 times (syndrom bits 0 1 2 3 4)
function [7-1:0] extended_hamming_code_43_36_f;
    input [36-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35];//16 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31]^in[34]^in[35];//16 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[35];//16 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28]^in[32]^in[33]^in[35];//16 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[35];//16 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33];//15 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32];//15 inputs
        extended_hamming_code_43_36_f = syndrom;
    end
endfunction
wire [7-1:0] stored_data_edc = extended_hamming_code_43_36_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_36_min_width (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [36-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_43_36_f
//Compute 7 bits Error Detection Code from a 36 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 8796093022208 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx   xx (16 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x  xx (16 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx   xx x (16 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx   xx x (16 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx   xx (16 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x x   (15 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xxx    (15 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
//  input bit 32 used 3 times (syndrom bits 2 3 6)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 1 4)
//  input bit 35 used 5 times (syndrom bits 0 1 2 3 4)
function [7-1:0] extended_hamming_code_43_36_f;
    input [36-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35];//16 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31]^in[34]^in[35];//16 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[35];//16 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28]^in[32]^in[33]^in[35];//16 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[35];//16 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33];//15 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32];//15 inputs
        extended_hamming_code_43_36_f = syndrom;
    end
endfunction
function [2+36-1:0] extended_hamming_code_43_36_f_correction_pattern_f;
    input [7-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [36-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {36{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			7'b0000000: begin
				correctable_error = 1'b0;
				correction_pattern = {36{1'b0}};
			end	
			7'b0000111: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 0]=1'b1;
			end
			7'b0111000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 1]=1'b1;
			end
			7'b1011000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 2]=1'b1;
			end
			7'b1100001: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 3]=1'b1;
			end
			7'b1000110: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 4]=1'b1;
			end
			7'b0100110: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 5]=1'b1;
			end
			7'b0011001: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 6]=1'b1;
			end
			7'b0001011: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 7]=1'b1;
			end
			7'b0110100: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 8]=1'b1;
			end
			7'b1010100: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 9]=1'b1;
			end
			7'b1101000: begin
				correction_pattern = {36{1'b0}};correction_pattern[10]=1'b1;
			end
			7'b1000011: begin
				correction_pattern = {36{1'b0}};correction_pattern[11]=1'b1;
			end
			7'b0100011: begin
				correction_pattern = {36{1'b0}};correction_pattern[12]=1'b1;
			end
			7'b0011100: begin
				correction_pattern = {36{1'b0}};correction_pattern[13]=1'b1;
			end
			7'b0011010: begin
				correction_pattern = {36{1'b0}};correction_pattern[14]=1'b1;
			end
			7'b0100101: begin
				correction_pattern = {36{1'b0}};correction_pattern[15]=1'b1;
			end
			7'b1000101: begin
				correction_pattern = {36{1'b0}};correction_pattern[16]=1'b1;
			end
			7'b1110000: begin
				correction_pattern = {36{1'b0}};correction_pattern[17]=1'b1;
			end
			7'b1001010: begin
				correction_pattern = {36{1'b0}};correction_pattern[18]=1'b1;
			end
			7'b0101010: begin
				correction_pattern = {36{1'b0}};correction_pattern[19]=1'b1;
			end
			7'b0010101: begin
				correction_pattern = {36{1'b0}};correction_pattern[20]=1'b1;
			end
			7'b0010110: begin
				correction_pattern = {36{1'b0}};correction_pattern[21]=1'b1;
			end
			7'b0101001: begin
				correction_pattern = {36{1'b0}};correction_pattern[22]=1'b1;
			end
			7'b1001001: begin
				correction_pattern = {36{1'b0}};correction_pattern[23]=1'b1;
			end
			7'b1100100: begin
				correction_pattern = {36{1'b0}};correction_pattern[24]=1'b1;
			end
			7'b1010010: begin
				correction_pattern = {36{1'b0}};correction_pattern[25]=1'b1;
			end
			7'b0110010: begin
				correction_pattern = {36{1'b0}};correction_pattern[26]=1'b1;
			end
			7'b0001101: begin
				correction_pattern = {36{1'b0}};correction_pattern[27]=1'b1;
			end
			7'b0001110: begin
				correction_pattern = {36{1'b0}};correction_pattern[28]=1'b1;
			end
			7'b0110001: begin
				correction_pattern = {36{1'b0}};correction_pattern[29]=1'b1;
			end
			7'b1010001: begin
				correction_pattern = {36{1'b0}};correction_pattern[30]=1'b1;
			end
			7'b1100010: begin
				correction_pattern = {36{1'b0}};correction_pattern[31]=1'b1;
			end
			7'b1001100: begin
				correction_pattern = {36{1'b0}};correction_pattern[32]=1'b1;
			end
			7'b0101100: begin
				correction_pattern = {36{1'b0}};correction_pattern[33]=1'b1;
			end
			7'b0010011: begin
				correction_pattern = {36{1'b0}};correction_pattern[34]=1'b1;
			end
			7'b0011111: begin
				correction_pattern = {36{1'b0}};correction_pattern[35]=1'b1;
			end
			7'b0000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b1000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_43_36_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [7-1:0] stored_data_edc = extended_hamming_code_43_36_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [36-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_43_36_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_40_min_width (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_46_40_f
//Compute 6 bits Error Detection Code from a 40 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 70368744177664 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[0]: x    x  xx x    x xx x  x xx  x xx x x x (18 inputs)
//  syndrom[1]: x     xx  x  x  xx x  x xx  xx  x xxx x  (18 inputs)
//  syndrom[2]:  x x    x x x   xx  xx x  x xx x x  xxxx (19 inputs)
//  syndrom[3]:  x  x x    x  xx x  x xx x x  x xx  xxxx (19 inputs)
//  syndrom[4]:   xx   x x    xx  xx  xx  xx x x  xx xx  (18 inputs)
//  syndrom[5]:   x xx      xx x  x xx  xx  x xx  xxx  x (18 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 2 4)
//  input bit  4 used 2 times (syndrom bits 3 5)
//  input bit  5 used 2 times (syndrom bits 0 5)
//  input bit  6 used 2 times (syndrom bits 1 3)
//  input bit  7 used 2 times (syndrom bits 1 4)
//  input bit  8 used 2 times (syndrom bits 0 2)
//  input bit  9 used 2 times (syndrom bits 0 4)
//  input bit 10 used 2 times (syndrom bits 1 2)
//  input bit 11 used 2 times (syndrom bits 0 3)
//  input bit 12 used 2 times (syndrom bits 2 5)
//  input bit 13 used 2 times (syndrom bits 1 5)
//  input bit 14 used 2 times (syndrom bits 3 4)
//  input bit 15 used 3 times (syndrom bits 3 4 5)
//  input bit 16 used 3 times (syndrom bits 0 1 2)
//  input bit 17 used 3 times (syndrom bits 1 2 3)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 0 1 4)
//  input bit 20 used 3 times (syndrom bits 2 3 5)
//  input bit 21 used 3 times (syndrom bits 0 2 5)
//  input bit 22 used 3 times (syndrom bits 1 3 4)
//  input bit 23 used 3 times (syndrom bits 2 3 4)
//  input bit 24 used 3 times (syndrom bits 0 1 5)
//  input bit 25 used 3 times (syndrom bits 1 3 5)
//  input bit 26 used 3 times (syndrom bits 0 2 4)
//  input bit 27 used 3 times (syndrom bits 0 3 4)
//  input bit 28 used 3 times (syndrom bits 1 2 5)
//  input bit 29 used 3 times (syndrom bits 1 2 4)
//  input bit 30 used 3 times (syndrom bits 0 3 5)
//  input bit 31 used 3 times (syndrom bits 2 4 5)
//  input bit 32 used 3 times (syndrom bits 0 1 3)
//  input bit 33 used 3 times (syndrom bits 0 2 3)
//  input bit 34 used 3 times (syndrom bits 1 4 5)
//  input bit 35 used 4 times (syndrom bits 0 1 4 5)
//  input bit 36 used 4 times (syndrom bits 1 2 3 5)
//  input bit 37 used 4 times (syndrom bits 0 2 3 4)
//  input bit 38 used 4 times (syndrom bits 1 2 3 4)
//  input bit 39 used 4 times (syndrom bits 0 2 3 5)
function [6-1:0] hamming_code_46_40_f;
    input [40-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 5]^in[ 8]^in[ 9]^in[11]^in[16]^in[18]^in[19]^in[21]^in[24]^in[26]^in[27]^in[30]^in[32]^in[33]^in[35]^in[37]^in[39];//18 inputs
        syndrom[1] = in[ 0]^in[ 6]^in[ 7]^in[10]^in[13]^in[16]^in[17]^in[19]^in[22]^in[24]^in[25]^in[28]^in[29]^in[32]^in[34]^in[35]^in[36]^in[38];//18 inputs
        syndrom[2] = in[ 1]^in[ 3]^in[ 8]^in[10]^in[12]^in[16]^in[17]^in[20]^in[21]^in[23]^in[26]^in[28]^in[29]^in[31]^in[33]^in[36]^in[37]^in[38]^in[39];//19 inputs
        syndrom[3] = in[ 1]^in[ 4]^in[ 6]^in[11]^in[14]^in[15]^in[17]^in[20]^in[22]^in[23]^in[25]^in[27]^in[30]^in[32]^in[33]^in[36]^in[37]^in[38]^in[39];//19 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 7]^in[ 9]^in[14]^in[15]^in[18]^in[19]^in[22]^in[23]^in[26]^in[27]^in[29]^in[31]^in[34]^in[35]^in[37]^in[38];//18 inputs
        syndrom[5] = in[ 2]^in[ 4]^in[ 5]^in[12]^in[13]^in[15]^in[18]^in[20]^in[21]^in[24]^in[25]^in[28]^in[30]^in[31]^in[34]^in[35]^in[36]^in[39];//18 inputs
        hamming_code_46_40_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = hamming_code_46_40_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_40_min_width (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_47_40_f
//Compute 7 bits Error Detection Code from a 40 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 140737488355328 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx   xxx x  (18 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x  xxxx   (18 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx   xx x xxx (19 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx   xx x xxx (19 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx   xxx  x (18 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x x  xxxx (19 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xxx   xxxx (19 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
//  input bit 32 used 3 times (syndrom bits 2 3 6)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 1 4)
//  input bit 35 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 36 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 37 used 5 times (syndrom bits 1 2 3 5 6)
//  input bit 38 used 5 times (syndrom bits 0 2 3 5 6)
//  input bit 39 used 5 times (syndrom bits 2 3 4 5 6)
function [7-1:0] extended_hamming_code_47_40_f;
    input [40-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35]^in[36]^in[38];//18 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31]^in[34]^in[35]^in[36]^in[37];//18 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39];//19 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39];//19 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[35]^in[36]^in[39];//18 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33]^in[36]^in[37]^in[38]^in[39];//19 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32]^in[36]^in[37]^in[38]^in[39];//19 inputs
        extended_hamming_code_47_40_f = syndrom;
    end
endfunction
wire [7-1:0] stored_data_edc = extended_hamming_code_47_40_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_40_min_width (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [40-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_47_40_f
//Compute 7 bits Error Detection Code from a 40 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 140737488355328 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx   xxx x  (18 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x  xxxx   (18 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx   xx x xxx (19 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx   xx x xxx (19 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx   xxx  x (18 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x x  xxxx (19 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xxx   xxxx (19 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
//  input bit 32 used 3 times (syndrom bits 2 3 6)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 1 4)
//  input bit 35 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 36 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 37 used 5 times (syndrom bits 1 2 3 5 6)
//  input bit 38 used 5 times (syndrom bits 0 2 3 5 6)
//  input bit 39 used 5 times (syndrom bits 2 3 4 5 6)
function [7-1:0] extended_hamming_code_47_40_f;
    input [40-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35]^in[36]^in[38];//18 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31]^in[34]^in[35]^in[36]^in[37];//18 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39];//19 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39];//19 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[35]^in[36]^in[39];//18 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33]^in[36]^in[37]^in[38]^in[39];//19 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32]^in[36]^in[37]^in[38]^in[39];//19 inputs
        extended_hamming_code_47_40_f = syndrom;
    end
endfunction
function [2+40-1:0] extended_hamming_code_47_40_f_correction_pattern_f;
    input [7-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [40-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {40{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			7'b0000000: begin
				correctable_error = 1'b0;
				correction_pattern = {40{1'b0}};
			end	
			7'b0000111: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 0]=1'b1;
			end
			7'b0111000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 1]=1'b1;
			end
			7'b1011000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 2]=1'b1;
			end
			7'b1100001: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 3]=1'b1;
			end
			7'b1000110: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 4]=1'b1;
			end
			7'b0100110: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 5]=1'b1;
			end
			7'b0011001: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 6]=1'b1;
			end
			7'b0001011: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 7]=1'b1;
			end
			7'b0110100: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 8]=1'b1;
			end
			7'b1010100: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 9]=1'b1;
			end
			7'b1101000: begin
				correction_pattern = {40{1'b0}};correction_pattern[10]=1'b1;
			end
			7'b1000011: begin
				correction_pattern = {40{1'b0}};correction_pattern[11]=1'b1;
			end
			7'b0100011: begin
				correction_pattern = {40{1'b0}};correction_pattern[12]=1'b1;
			end
			7'b0011100: begin
				correction_pattern = {40{1'b0}};correction_pattern[13]=1'b1;
			end
			7'b0011010: begin
				correction_pattern = {40{1'b0}};correction_pattern[14]=1'b1;
			end
			7'b0100101: begin
				correction_pattern = {40{1'b0}};correction_pattern[15]=1'b1;
			end
			7'b1000101: begin
				correction_pattern = {40{1'b0}};correction_pattern[16]=1'b1;
			end
			7'b1110000: begin
				correction_pattern = {40{1'b0}};correction_pattern[17]=1'b1;
			end
			7'b1001010: begin
				correction_pattern = {40{1'b0}};correction_pattern[18]=1'b1;
			end
			7'b0101010: begin
				correction_pattern = {40{1'b0}};correction_pattern[19]=1'b1;
			end
			7'b0010101: begin
				correction_pattern = {40{1'b0}};correction_pattern[20]=1'b1;
			end
			7'b0010110: begin
				correction_pattern = {40{1'b0}};correction_pattern[21]=1'b1;
			end
			7'b0101001: begin
				correction_pattern = {40{1'b0}};correction_pattern[22]=1'b1;
			end
			7'b1001001: begin
				correction_pattern = {40{1'b0}};correction_pattern[23]=1'b1;
			end
			7'b1100100: begin
				correction_pattern = {40{1'b0}};correction_pattern[24]=1'b1;
			end
			7'b1010010: begin
				correction_pattern = {40{1'b0}};correction_pattern[25]=1'b1;
			end
			7'b0110010: begin
				correction_pattern = {40{1'b0}};correction_pattern[26]=1'b1;
			end
			7'b0001101: begin
				correction_pattern = {40{1'b0}};correction_pattern[27]=1'b1;
			end
			7'b0001110: begin
				correction_pattern = {40{1'b0}};correction_pattern[28]=1'b1;
			end
			7'b0110001: begin
				correction_pattern = {40{1'b0}};correction_pattern[29]=1'b1;
			end
			7'b1010001: begin
				correction_pattern = {40{1'b0}};correction_pattern[30]=1'b1;
			end
			7'b1100010: begin
				correction_pattern = {40{1'b0}};correction_pattern[31]=1'b1;
			end
			7'b1001100: begin
				correction_pattern = {40{1'b0}};correction_pattern[32]=1'b1;
			end
			7'b0101100: begin
				correction_pattern = {40{1'b0}};correction_pattern[33]=1'b1;
			end
			7'b0010011: begin
				correction_pattern = {40{1'b0}};correction_pattern[34]=1'b1;
			end
			7'b0011111: begin
				correction_pattern = {40{1'b0}};correction_pattern[35]=1'b1;
			end
			7'b1110011: begin
				correction_pattern = {40{1'b0}};correction_pattern[36]=1'b1;
			end
			7'b1101110: begin
				correction_pattern = {40{1'b0}};correction_pattern[37]=1'b1;
			end
			7'b1101101: begin
				correction_pattern = {40{1'b0}};correction_pattern[38]=1'b1;
			end
			7'b1111100: begin
				correction_pattern = {40{1'b0}};correction_pattern[39]=1'b1;
			end
			7'b0000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b1000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_47_40_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [7-1:0] stored_data_edc = extended_hamming_code_47_40_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [40-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_47_40_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_48_min_width (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_54_48_f
//Compute 6 bits Error Detection Code from a 48 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 18014398509481984 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[0]: x    x  xx x    x xx x  x xx  x xx x x xxxx  xxx (24 inputs)
//  syndrom[1]: x     xx  x  x  xx x  x xx  xx  x x x x  xxxxxxx (24 inputs)
//  syndrom[2]:  x x    x x x   xx  xx x  x xx x x xxxxx xx x  x (24 inputs)
//  syndrom[3]:  x  x x    x  xx x  x xx x x  x xx  xxxxx  x xxx (24 inputs)
//  syndrom[4]:   xx   x x    xx  xx  xx  xx x x  xx xx x xxxx   (23 inputs)
//  syndrom[5]:   x xx      xx x  x xx  xx  x xx  xxx  xxx xx x  (23 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 2 4)
//  input bit  4 used 2 times (syndrom bits 3 5)
//  input bit  5 used 2 times (syndrom bits 0 5)
//  input bit  6 used 2 times (syndrom bits 1 3)
//  input bit  7 used 2 times (syndrom bits 1 4)
//  input bit  8 used 2 times (syndrom bits 0 2)
//  input bit  9 used 2 times (syndrom bits 0 4)
//  input bit 10 used 2 times (syndrom bits 1 2)
//  input bit 11 used 2 times (syndrom bits 0 3)
//  input bit 12 used 2 times (syndrom bits 2 5)
//  input bit 13 used 2 times (syndrom bits 1 5)
//  input bit 14 used 2 times (syndrom bits 3 4)
//  input bit 15 used 3 times (syndrom bits 3 4 5)
//  input bit 16 used 3 times (syndrom bits 0 1 2)
//  input bit 17 used 3 times (syndrom bits 1 2 3)
//  input bit 18 used 3 times (syndrom bits 0 4 5)
//  input bit 19 used 3 times (syndrom bits 0 1 4)
//  input bit 20 used 3 times (syndrom bits 2 3 5)
//  input bit 21 used 3 times (syndrom bits 0 2 5)
//  input bit 22 used 3 times (syndrom bits 1 3 4)
//  input bit 23 used 3 times (syndrom bits 2 3 4)
//  input bit 24 used 3 times (syndrom bits 0 1 5)
//  input bit 25 used 3 times (syndrom bits 1 3 5)
//  input bit 26 used 3 times (syndrom bits 0 2 4)
//  input bit 27 used 3 times (syndrom bits 0 3 4)
//  input bit 28 used 3 times (syndrom bits 1 2 5)
//  input bit 29 used 3 times (syndrom bits 1 2 4)
//  input bit 30 used 3 times (syndrom bits 0 3 5)
//  input bit 31 used 3 times (syndrom bits 2 4 5)
//  input bit 32 used 3 times (syndrom bits 0 1 3)
//  input bit 33 used 3 times (syndrom bits 0 2 3)
//  input bit 34 used 3 times (syndrom bits 1 4 5)
//  input bit 35 used 4 times (syndrom bits 0 2 4 5)
//  input bit 36 used 4 times (syndrom bits 1 2 3 5)
//  input bit 37 used 4 times (syndrom bits 0 2 3 4)
//  input bit 38 used 4 times (syndrom bits 1 2 3 4)
//  input bit 39 used 4 times (syndrom bits 0 2 3 5)
//  input bit 40 used 4 times (syndrom bits 0 3 4 5)
//  input bit 41 used 4 times (syndrom bits 0 1 2 5)
//  input bit 42 used 4 times (syndrom bits 0 1 2 4)
//  input bit 43 used 4 times (syndrom bits 1 3 4 5)
//  input bit 44 used 4 times (syndrom bits 1 2 4 5)
//  input bit 45 used 4 times (syndrom bits 0 1 3 4)
//  input bit 46 used 4 times (syndrom bits 0 1 3 5)
//  input bit 47 used 4 times (syndrom bits 0 1 2 3)
function [6-1:0] hamming_code_54_48_f;
    input [48-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 5]^in[ 8]^in[ 9]^in[11]^in[16]^in[18]^in[19]^in[21]^in[24]^in[26]^in[27]^in[30]^in[32]^in[33]^in[35]^in[37]^in[39]^in[40]^in[41]^in[42]^in[45]^in[46]^in[47];//24 inputs
        syndrom[1] = in[ 0]^in[ 6]^in[ 7]^in[10]^in[13]^in[16]^in[17]^in[19]^in[22]^in[24]^in[25]^in[28]^in[29]^in[32]^in[34]^in[36]^in[38]^in[41]^in[42]^in[43]^in[44]^in[45]^in[46]^in[47];//24 inputs
        syndrom[2] = in[ 1]^in[ 3]^in[ 8]^in[10]^in[12]^in[16]^in[17]^in[20]^in[21]^in[23]^in[26]^in[28]^in[29]^in[31]^in[33]^in[35]^in[36]^in[37]^in[38]^in[39]^in[41]^in[42]^in[44]^in[47];//24 inputs
        syndrom[3] = in[ 1]^in[ 4]^in[ 6]^in[11]^in[14]^in[15]^in[17]^in[20]^in[22]^in[23]^in[25]^in[27]^in[30]^in[32]^in[33]^in[36]^in[37]^in[38]^in[39]^in[40]^in[43]^in[45]^in[46]^in[47];//24 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 7]^in[ 9]^in[14]^in[15]^in[18]^in[19]^in[22]^in[23]^in[26]^in[27]^in[29]^in[31]^in[34]^in[35]^in[37]^in[38]^in[40]^in[42]^in[43]^in[44]^in[45];//23 inputs
        syndrom[5] = in[ 2]^in[ 4]^in[ 5]^in[12]^in[13]^in[15]^in[18]^in[20]^in[21]^in[24]^in[25]^in[28]^in[30]^in[31]^in[34]^in[35]^in[36]^in[39]^in[40]^in[41]^in[43]^in[44]^in[46];//23 inputs
        hamming_code_54_48_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = hamming_code_54_48_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_48_min_width (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_55_48_f
//Compute 7 bits Error Detection Code from a 48 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 36028797018963968 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx   xxx x xxxxx xx (25 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x  xxxx  xxxx xxx (25 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx   xx x xxxx x  xxx (24 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx   xx x xxx x xxxx  (24 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx   xxx  xxxxxxx   (24 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x x  xxxxx  xxx x (24 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xxx   xxxx xx x xx (24 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
//  input bit 32 used 3 times (syndrom bits 2 3 6)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 1 4)
//  input bit 35 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 36 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 37 used 5 times (syndrom bits 1 2 3 5 6)
//  input bit 38 used 5 times (syndrom bits 0 2 3 5 6)
//  input bit 39 used 5 times (syndrom bits 2 3 4 5 6)
//  input bit 40 used 5 times (syndrom bits 0 1 2 4 5)
//  input bit 41 used 5 times (syndrom bits 0 1 3 4 6)
//  input bit 42 used 5 times (syndrom bits 0 1 2 4 6)
//  input bit 43 used 5 times (syndrom bits 0 1 3 4 5)
//  input bit 44 used 5 times (syndrom bits 0 3 4 5 6)
//  input bit 45 used 5 times (syndrom bits 1 2 3 4 5)
//  input bit 46 used 5 times (syndrom bits 0 1 2 3 6)
//  input bit 47 used 5 times (syndrom bits 0 1 2 5 6)
function [7-1:0] extended_hamming_code_55_48_f;
    input [48-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35]^in[36]^in[38]^in[40]^in[41]^in[42]^in[43]^in[44]^in[46]^in[47];//25 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31]^in[34]^in[35]^in[36]^in[37]^in[40]^in[41]^in[42]^in[43]^in[45]^in[46]^in[47];//25 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39]^in[40]^in[42]^in[45]^in[46]^in[47];//24 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39]^in[41]^in[43]^in[44]^in[45]^in[46];//24 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[35]^in[36]^in[39]^in[40]^in[41]^in[42]^in[43]^in[44]^in[45];//24 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33]^in[36]^in[37]^in[38]^in[39]^in[40]^in[43]^in[44]^in[45]^in[47];//24 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32]^in[36]^in[37]^in[38]^in[39]^in[41]^in[42]^in[44]^in[46]^in[47];//24 inputs
        extended_hamming_code_55_48_f = syndrom;
    end
endfunction
wire [7-1:0] stored_data_edc = extended_hamming_code_55_48_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_48_min_width (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [48-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_55_48_f
//Compute 7 bits Error Detection Code from a 48 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 36028797018963968 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[0]: x  x  xx   xx  xx   x xx   x xx   xxx x xxxxx xx (25 inputs)
//  syndrom[1]: x   xx x   xx x   xx x   xx x  x  xxxx  xxxx xxx (25 inputs)
//  syndrom[2]: x   xx  xx   x xx   xx  x  xx   xx x xxxx x  xxx (24 inputs)
//  syndrom[3]:  xx   xx  x  xx   xx  xx   xx   xx x xxx x xxxx  (24 inputs)
//  syndrom[4]:  xx   x xx   xx  x  xx   xx  xx   xxx  xxxxxxx   (24 inputs)
//  syndrom[5]:  x x x  x x x  x x x  x x x  x x x  xxxxx  xxx x (24 inputs)
//  syndrom[6]:   xxx    xxx    xxx    xxx    xxx   xxxx xx x xx (24 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 4 6)
//  input bit  3 used 3 times (syndrom bits 0 5 6)
//  input bit  4 used 3 times (syndrom bits 1 2 6)
//  input bit  5 used 3 times (syndrom bits 1 2 5)
//  input bit  6 used 3 times (syndrom bits 0 3 4)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 2 4 5)
//  input bit  9 used 3 times (syndrom bits 2 4 6)
//  input bit 10 used 3 times (syndrom bits 3 5 6)
//  input bit 11 used 3 times (syndrom bits 0 1 6)
//  input bit 12 used 3 times (syndrom bits 0 1 5)
//  input bit 13 used 3 times (syndrom bits 2 3 4)
//  input bit 14 used 3 times (syndrom bits 1 3 4)
//  input bit 15 used 3 times (syndrom bits 0 2 5)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 4 5 6)
//  input bit 18 used 3 times (syndrom bits 1 3 6)
//  input bit 19 used 3 times (syndrom bits 1 3 5)
//  input bit 20 used 3 times (syndrom bits 0 2 4)
//  input bit 21 used 3 times (syndrom bits 1 2 4)
//  input bit 22 used 3 times (syndrom bits 0 3 5)
//  input bit 23 used 3 times (syndrom bits 0 3 6)
//  input bit 24 used 3 times (syndrom bits 2 5 6)
//  input bit 25 used 3 times (syndrom bits 1 4 6)
//  input bit 26 used 3 times (syndrom bits 1 4 5)
//  input bit 27 used 3 times (syndrom bits 0 2 3)
//  input bit 28 used 3 times (syndrom bits 1 2 3)
//  input bit 29 used 3 times (syndrom bits 0 4 5)
//  input bit 30 used 3 times (syndrom bits 0 4 6)
//  input bit 31 used 3 times (syndrom bits 1 5 6)
//  input bit 32 used 3 times (syndrom bits 2 3 6)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 1 4)
//  input bit 35 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 36 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 37 used 5 times (syndrom bits 1 2 3 5 6)
//  input bit 38 used 5 times (syndrom bits 0 2 3 5 6)
//  input bit 39 used 5 times (syndrom bits 2 3 4 5 6)
//  input bit 40 used 5 times (syndrom bits 0 1 2 4 5)
//  input bit 41 used 5 times (syndrom bits 0 1 3 4 6)
//  input bit 42 used 5 times (syndrom bits 0 1 2 4 6)
//  input bit 43 used 5 times (syndrom bits 0 1 3 4 5)
//  input bit 44 used 5 times (syndrom bits 0 3 4 5 6)
//  input bit 45 used 5 times (syndrom bits 1 2 3 4 5)
//  input bit 46 used 5 times (syndrom bits 0 1 2 3 6)
//  input bit 47 used 5 times (syndrom bits 0 1 2 5 6)
function [7-1:0] extended_hamming_code_55_48_f;
    input [48-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 3]^in[ 6]^in[ 7]^in[11]^in[12]^in[15]^in[16]^in[20]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35]^in[36]^in[38]^in[40]^in[41]^in[42]^in[43]^in[44]^in[46]^in[47];//25 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 5]^in[ 7]^in[11]^in[12]^in[14]^in[18]^in[19]^in[21]^in[25]^in[26]^in[28]^in[31]^in[34]^in[35]^in[36]^in[37]^in[40]^in[41]^in[42]^in[43]^in[45]^in[46]^in[47];//25 inputs
        syndrom[2] = in[ 0]^in[ 4]^in[ 5]^in[ 8]^in[ 9]^in[13]^in[15]^in[16]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39]^in[40]^in[42]^in[45]^in[46]^in[47];//24 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 6]^in[ 7]^in[10]^in[13]^in[14]^in[18]^in[19]^in[22]^in[23]^in[27]^in[28]^in[32]^in[33]^in[35]^in[37]^in[38]^in[39]^in[41]^in[43]^in[44]^in[45]^in[46];//24 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 6]^in[ 8]^in[ 9]^in[13]^in[14]^in[17]^in[20]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[35]^in[36]^in[39]^in[40]^in[41]^in[42]^in[43]^in[44]^in[45];//24 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 5]^in[ 8]^in[10]^in[12]^in[15]^in[17]^in[19]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33]^in[36]^in[37]^in[38]^in[39]^in[40]^in[43]^in[44]^in[45]^in[47];//24 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 4]^in[ 9]^in[10]^in[11]^in[16]^in[17]^in[18]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32]^in[36]^in[37]^in[38]^in[39]^in[41]^in[42]^in[44]^in[46]^in[47];//24 inputs
        extended_hamming_code_55_48_f = syndrom;
    end
endfunction
function [2+48-1:0] extended_hamming_code_55_48_f_correction_pattern_f;
    input [7-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [48-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {48{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			7'b0000000: begin
				correctable_error = 1'b0;
				correction_pattern = {48{1'b0}};
			end	
			7'b0000111: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 0]=1'b1;
			end
			7'b0111000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 1]=1'b1;
			end
			7'b1011000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 2]=1'b1;
			end
			7'b1100001: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 3]=1'b1;
			end
			7'b1000110: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 4]=1'b1;
			end
			7'b0100110: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 5]=1'b1;
			end
			7'b0011001: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 6]=1'b1;
			end
			7'b0001011: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 7]=1'b1;
			end
			7'b0110100: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 8]=1'b1;
			end
			7'b1010100: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 9]=1'b1;
			end
			7'b1101000: begin
				correction_pattern = {48{1'b0}};correction_pattern[10]=1'b1;
			end
			7'b1000011: begin
				correction_pattern = {48{1'b0}};correction_pattern[11]=1'b1;
			end
			7'b0100011: begin
				correction_pattern = {48{1'b0}};correction_pattern[12]=1'b1;
			end
			7'b0011100: begin
				correction_pattern = {48{1'b0}};correction_pattern[13]=1'b1;
			end
			7'b0011010: begin
				correction_pattern = {48{1'b0}};correction_pattern[14]=1'b1;
			end
			7'b0100101: begin
				correction_pattern = {48{1'b0}};correction_pattern[15]=1'b1;
			end
			7'b1000101: begin
				correction_pattern = {48{1'b0}};correction_pattern[16]=1'b1;
			end
			7'b1110000: begin
				correction_pattern = {48{1'b0}};correction_pattern[17]=1'b1;
			end
			7'b1001010: begin
				correction_pattern = {48{1'b0}};correction_pattern[18]=1'b1;
			end
			7'b0101010: begin
				correction_pattern = {48{1'b0}};correction_pattern[19]=1'b1;
			end
			7'b0010101: begin
				correction_pattern = {48{1'b0}};correction_pattern[20]=1'b1;
			end
			7'b0010110: begin
				correction_pattern = {48{1'b0}};correction_pattern[21]=1'b1;
			end
			7'b0101001: begin
				correction_pattern = {48{1'b0}};correction_pattern[22]=1'b1;
			end
			7'b1001001: begin
				correction_pattern = {48{1'b0}};correction_pattern[23]=1'b1;
			end
			7'b1100100: begin
				correction_pattern = {48{1'b0}};correction_pattern[24]=1'b1;
			end
			7'b1010010: begin
				correction_pattern = {48{1'b0}};correction_pattern[25]=1'b1;
			end
			7'b0110010: begin
				correction_pattern = {48{1'b0}};correction_pattern[26]=1'b1;
			end
			7'b0001101: begin
				correction_pattern = {48{1'b0}};correction_pattern[27]=1'b1;
			end
			7'b0001110: begin
				correction_pattern = {48{1'b0}};correction_pattern[28]=1'b1;
			end
			7'b0110001: begin
				correction_pattern = {48{1'b0}};correction_pattern[29]=1'b1;
			end
			7'b1010001: begin
				correction_pattern = {48{1'b0}};correction_pattern[30]=1'b1;
			end
			7'b1100010: begin
				correction_pattern = {48{1'b0}};correction_pattern[31]=1'b1;
			end
			7'b1001100: begin
				correction_pattern = {48{1'b0}};correction_pattern[32]=1'b1;
			end
			7'b0101100: begin
				correction_pattern = {48{1'b0}};correction_pattern[33]=1'b1;
			end
			7'b0010011: begin
				correction_pattern = {48{1'b0}};correction_pattern[34]=1'b1;
			end
			7'b0011111: begin
				correction_pattern = {48{1'b0}};correction_pattern[35]=1'b1;
			end
			7'b1110011: begin
				correction_pattern = {48{1'b0}};correction_pattern[36]=1'b1;
			end
			7'b1101110: begin
				correction_pattern = {48{1'b0}};correction_pattern[37]=1'b1;
			end
			7'b1101101: begin
				correction_pattern = {48{1'b0}};correction_pattern[38]=1'b1;
			end
			7'b1111100: begin
				correction_pattern = {48{1'b0}};correction_pattern[39]=1'b1;
			end
			7'b0110111: begin
				correction_pattern = {48{1'b0}};correction_pattern[40]=1'b1;
			end
			7'b1011011: begin
				correction_pattern = {48{1'b0}};correction_pattern[41]=1'b1;
			end
			7'b1010111: begin
				correction_pattern = {48{1'b0}};correction_pattern[42]=1'b1;
			end
			7'b0111011: begin
				correction_pattern = {48{1'b0}};correction_pattern[43]=1'b1;
			end
			7'b1111001: begin
				correction_pattern = {48{1'b0}};correction_pattern[44]=1'b1;
			end
			7'b0111110: begin
				correction_pattern = {48{1'b0}};correction_pattern[45]=1'b1;
			end
			7'b1001111: begin
				correction_pattern = {48{1'b0}};correction_pattern[46]=1'b1;
			end
			7'b1100111: begin
				correction_pattern = {48{1'b0}};correction_pattern[47]=1'b1;
			end
			7'b0000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b0100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			7'b1000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_55_48_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [7-1:0] stored_data_edc = extended_hamming_code_55_48_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [48-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_55_48_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_64_min_width (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_71_64_f
//Compute 7 bits Error Detection Code from a 64 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 2361183241434822606848 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[0]: x    x x    xx      xx   xx x   xx x   xx x   xx x  x  xxx   xxx (26 inputs)
//  syndrom[1]: x     x xx      xx     xxx    xxx    xxx    xxx    xxx   xx xx   (25 inputs)
//  syndrom[2]:  x   x  x x    x  x   x x x  x x x  x x x  x x x  x x x  xxx  x  (25 inputs)
//  syndrom[3]:  x    xx   x  x    x  xx   xx  x  xx   xx  xx   xx   xx  xxx  xx (26 inputs)
//  syndrom[4]:   xx       xx    xx   xx   x xx   xx  x  xx   xx  xx   xx  xxx x (26 inputs)
//  syndrom[5]:   x x     x  x  x  x x   xx  xx   x xx   xx  x  xx   xx x  xxx   (25 inputs)
//  syndrom[6]:    xx    x    xx    xx  x  xx   xx  xx   x xx   x xx   xx x x xx (26 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 4 6)
//  input bit  4 used 2 times (syndrom bits 5 6)
//  input bit  5 used 2 times (syndrom bits 0 2)
//  input bit  6 used 2 times (syndrom bits 1 3)
//  input bit  7 used 2 times (syndrom bits 0 3)
//  input bit  8 used 2 times (syndrom bits 1 2)
//  input bit  9 used 2 times (syndrom bits 1 6)
//  input bit 10 used 2 times (syndrom bits 2 5)
//  input bit 11 used 2 times (syndrom bits 3 4)
//  input bit 12 used 2 times (syndrom bits 0 4)
//  input bit 13 used 2 times (syndrom bits 0 5)
//  input bit 14 used 2 times (syndrom bits 3 6)
//  input bit 15 used 2 times (syndrom bits 2 6)
//  input bit 16 used 2 times (syndrom bits 1 5)
//  input bit 17 used 2 times (syndrom bits 1 4)
//  input bit 18 used 2 times (syndrom bits 2 4)
//  input bit 19 used 2 times (syndrom bits 3 5)
//  input bit 20 used 2 times (syndrom bits 0 6)
//  input bit 21 used 3 times (syndrom bits 0 5 6)
//  input bit 22 used 3 times (syndrom bits 2 3 4)
//  input bit 23 used 3 times (syndrom bits 1 3 4)
//  input bit 24 used 3 times (syndrom bits 1 2 6)
//  input bit 25 used 3 times (syndrom bits 0 1 5)
//  input bit 26 used 3 times (syndrom bits 0 2 5)
//  input bit 27 used 3 times (syndrom bits 3 4 6)
//  input bit 28 used 3 times (syndrom bits 0 3 6)
//  input bit 29 used 3 times (syndrom bits 2 4 5)
//  input bit 30 used 3 times (syndrom bits 1 4 5)
//  input bit 31 used 3 times (syndrom bits 1 2 3)
//  input bit 32 used 3 times (syndrom bits 0 1 6)
//  input bit 33 used 3 times (syndrom bits 0 2 6)
//  input bit 34 used 3 times (syndrom bits 3 4 5)
//  input bit 35 used 3 times (syndrom bits 0 3 4)
//  input bit 36 used 3 times (syndrom bits 2 5 6)
//  input bit 37 used 3 times (syndrom bits 1 5 6)
//  input bit 38 used 3 times (syndrom bits 1 2 4)
//  input bit 39 used 3 times (syndrom bits 0 1 3)
//  input bit 40 used 3 times (syndrom bits 0 2 3)
//  input bit 41 used 3 times (syndrom bits 4 5 6)
//  input bit 42 used 3 times (syndrom bits 0 4 5)
//  input bit 43 used 3 times (syndrom bits 2 3 6)
//  input bit 44 used 3 times (syndrom bits 1 3 6)
//  input bit 45 used 3 times (syndrom bits 1 2 5)
//  input bit 46 used 3 times (syndrom bits 0 1 4)
//  input bit 47 used 3 times (syndrom bits 0 2 4)
//  input bit 48 used 3 times (syndrom bits 3 5 6)
//  input bit 49 used 3 times (syndrom bits 0 3 5)
//  input bit 50 used 3 times (syndrom bits 2 4 6)
//  input bit 51 used 3 times (syndrom bits 1 4 6)
//  input bit 52 used 3 times (syndrom bits 0 1 2)
//  input bit 53 used 3 times (syndrom bits 1 3 5)
//  input bit 54 used 3 times (syndrom bits 2 3 5)
//  input bit 55 used 3 times (syndrom bits 0 4 6)
//  input bit 56 used 4 times (syndrom bits 0 4 5 6)
//  input bit 57 used 4 times (syndrom bits 0 1 2 3)
//  input bit 58 used 4 times (syndrom bits 1 2 3 6)
//  input bit 59 used 4 times (syndrom bits 2 3 4 5)
//  input bit 60 used 4 times (syndrom bits 1 4 5 6)
//  input bit 61 used 4 times (syndrom bits 0 1 4 5)
//  input bit 62 used 4 times (syndrom bits 0 2 3 6)
//  input bit 63 used 4 times (syndrom bits 0 3 4 6)
function [7-1:0] hamming_code_71_64_f;
    input [64-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 5]^in[ 7]^in[12]^in[13]^in[20]^in[21]^in[25]^in[26]^in[28]^in[32]^in[33]^in[35]^in[39]^in[40]^in[42]^in[46]^in[47]^in[49]^in[52]^in[55]^in[56]^in[57]^in[61]^in[62]^in[63];//26 inputs
        syndrom[1] = in[ 0]^in[ 6]^in[ 8]^in[ 9]^in[16]^in[17]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32]^in[37]^in[38]^in[39]^in[44]^in[45]^in[46]^in[51]^in[52]^in[53]^in[57]^in[58]^in[60]^in[61];//25 inputs
        syndrom[2] = in[ 1]^in[ 5]^in[ 8]^in[10]^in[15]^in[18]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33]^in[36]^in[38]^in[40]^in[43]^in[45]^in[47]^in[50]^in[52]^in[54]^in[57]^in[58]^in[59]^in[62];//25 inputs
        syndrom[3] = in[ 1]^in[ 6]^in[ 7]^in[11]^in[14]^in[19]^in[22]^in[23]^in[27]^in[28]^in[31]^in[34]^in[35]^in[39]^in[40]^in[43]^in[44]^in[48]^in[49]^in[53]^in[54]^in[57]^in[58]^in[59]^in[62]^in[63];//26 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[11]^in[12]^in[17]^in[18]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35]^in[38]^in[41]^in[42]^in[46]^in[47]^in[50]^in[51]^in[55]^in[56]^in[59]^in[60]^in[61]^in[63];//26 inputs
        syndrom[5] = in[ 2]^in[ 4]^in[10]^in[13]^in[16]^in[19]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[36]^in[37]^in[41]^in[42]^in[45]^in[48]^in[49]^in[53]^in[54]^in[56]^in[59]^in[60]^in[61];//25 inputs
        syndrom[6] = in[ 3]^in[ 4]^in[ 9]^in[14]^in[15]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[36]^in[37]^in[41]^in[43]^in[44]^in[48]^in[50]^in[51]^in[55]^in[56]^in[58]^in[60]^in[62]^in[63];//26 inputs
        hamming_code_71_64_f = syndrom;
    end
endfunction
wire [7-1:0] stored_data_edc = hamming_code_71_64_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_64_min_width (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_72_64_f
//Compute 8 bits Error Detection Code from a 64 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[0]: x   xx    xx   xx   x x  x  xx    xx  x x  x   x  xx  x x  xxxx  (26 inputs)
//  syndrom[1]: x   x x  x  xx   x  xx    xx   xx   x  xx    x xx    xx x x xxx  (26 inputs)
//  syndrom[2]: x    xx x    xx x    xx x    xx  x  xx    x x x   x xx   xxx x x (26 inputs)
//  syndrom[3]:  xx    x xx    x xx    x xx    x xx     xxx x     x xx   xxx  xx (26 inputs)
//  syndrom[4]:  x x   xx   x x  x x   xx   xx    xxx      xxx  xx    x  xxxx  x (26 inputs)
//  syndrom[5]:  x  xx    xx  x   xx x    xx  x  x x   x x   xx  x x   xxx  xx x (26 inputs)
//  syndrom[6]:   xx  x  x x   xx   x  xx   x x x    xxx x      xx  x  xxx  xxx  (26 inputs)
//  syndrom[7]:   xx   xx   xx    xx  x  x x   xx    xx   xx  xx   x   xx xx  xx (26 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 6 7)
//  input bit  3 used 3 times (syndrom bits 4 6 7)
//  input bit  4 used 3 times (syndrom bits 0 1 5)
//  input bit  5 used 3 times (syndrom bits 0 2 5)
//  input bit  6 used 3 times (syndrom bits 1 2 6)
//  input bit  7 used 3 times (syndrom bits 3 4 7)
//  input bit  8 used 3 times (syndrom bits 2 4 7)
//  input bit  9 used 3 times (syndrom bits 1 3 6)
//  input bit 10 used 3 times (syndrom bits 0 3 5)
//  input bit 11 used 3 times (syndrom bits 0 5 6)
//  input bit 12 used 3 times (syndrom bits 1 4 7)
//  input bit 13 used 3 times (syndrom bits 1 2 7)
//  input bit 14 used 3 times (syndrom bits 2 4 5)
//  input bit 15 used 3 times (syndrom bits 0 3 6)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 1 3 4)
//  input bit 18 used 3 times (syndrom bits 3 5 7)
//  input bit 19 used 3 times (syndrom bits 4 5 7)
//  input bit 20 used 3 times (syndrom bits 0 1 6)
//  input bit 21 used 3 times (syndrom bits 1 2 5)
//  input bit 22 used 3 times (syndrom bits 0 2 7)
//  input bit 23 used 3 times (syndrom bits 3 4 6)
//  input bit 24 used 3 times (syndrom bits 2 4 6)
//  input bit 25 used 3 times (syndrom bits 0 3 7)
//  input bit 26 used 3 times (syndrom bits 1 3 5)
//  input bit 27 used 3 times (syndrom bits 1 5 7)
//  input bit 28 used 3 times (syndrom bits 0 4 6)
//  input bit 29 used 3 times (syndrom bits 0 2 4)
//  input bit 30 used 3 times (syndrom bits 2 5 6)
//  input bit 31 used 3 times (syndrom bits 1 3 7)
//  input bit 32 used 3 times (syndrom bits 1 6 7)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 3 4)
//  input bit 35 used 3 times (syndrom bits 0 4 5)
//  input bit 36 used 3 times (syndrom bits 1 2 4)
//  input bit 37 used 3 times (syndrom bits 2 6 7)
//  input bit 38 used 3 times (syndrom bits 0 6 7)
//  input bit 39 used 3 times (syndrom bits 1 5 6)
//  input bit 40 used 3 times (syndrom bits 0 1 3)
//  input bit 41 used 3 times (syndrom bits 3 5 6)
//  input bit 42 used 3 times (syndrom bits 2 3 7)
//  input bit 43 used 3 times (syndrom bits 0 4 7)
//  input bit 44 used 3 times (syndrom bits 2 3 4)
//  input bit 45 used 3 times (syndrom bits 1 4 5)
//  input bit 46 used 3 times (syndrom bits 2 5 7)
//  input bit 47 used 3 times (syndrom bits 0 1 7)
//  input bit 48 used 3 times (syndrom bits 1 4 6)
//  input bit 49 used 3 times (syndrom bits 4 5 6)
//  input bit 50 used 3 times (syndrom bits 0 2 3)
//  input bit 51 used 3 times (syndrom bits 0 5 7)
//  input bit 52 used 3 times (syndrom bits 2 3 6)
//  input bit 53 used 3 times (syndrom bits 1 2 3)
//  input bit 54 used 3 times (syndrom bits 0 1 4)
//  input bit 55 used 3 times (syndrom bits 5 6 7)
//  input bit 56 used 5 times (syndrom bits 0 1 5 6 7)
//  input bit 57 used 5 times (syndrom bits 2 3 4 5 6)
//  input bit 58 used 5 times (syndrom bits 1 2 3 4 7)
//  input bit 59 used 5 times (syndrom bits 0 2 3 4 7)
//  input bit 60 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 61 used 5 times (syndrom bits 0 1 2 5 6)
//  input bit 62 used 5 times (syndrom bits 0 1 3 6 7)
//  input bit 63 used 5 times (syndrom bits 2 3 4 5 7)
function [8-1:0] extended_hamming_code_72_64_f;
    input [64-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 5]^in[10]^in[11]^in[15]^in[16]^in[20]^in[22]^in[25]^in[28]^in[29]^in[34]^in[35]^in[38]^in[40]^in[43]^in[47]^in[50]^in[51]^in[54]^in[56]^in[59]^in[60]^in[61]^in[62];//26 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 6]^in[ 9]^in[12]^in[13]^in[17]^in[20]^in[21]^in[26]^in[27]^in[31]^in[32]^in[36]^in[39]^in[40]^in[45]^in[47]^in[48]^in[53]^in[54]^in[56]^in[58]^in[60]^in[61]^in[62];//26 inputs
        syndrom[2] = in[ 0]^in[ 5]^in[ 6]^in[ 8]^in[13]^in[14]^in[16]^in[21]^in[22]^in[24]^in[29]^in[30]^in[33]^in[36]^in[37]^in[42]^in[44]^in[46]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[61]^in[63];//26 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 7]^in[ 9]^in[10]^in[15]^in[17]^in[18]^in[23]^in[25]^in[26]^in[31]^in[33]^in[34]^in[40]^in[41]^in[42]^in[44]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[62]^in[63];//26 inputs
        syndrom[4] = in[ 1]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[14]^in[17]^in[19]^in[23]^in[24]^in[28]^in[29]^in[34]^in[35]^in[36]^in[43]^in[44]^in[45]^in[48]^in[49]^in[54]^in[57]^in[58]^in[59]^in[60]^in[63];//26 inputs
        syndrom[5] = in[ 1]^in[ 4]^in[ 5]^in[10]^in[11]^in[14]^in[18]^in[19]^in[21]^in[26]^in[27]^in[30]^in[33]^in[35]^in[39]^in[41]^in[45]^in[46]^in[49]^in[51]^in[55]^in[56]^in[57]^in[60]^in[61]^in[63];//26 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 6]^in[ 9]^in[11]^in[15]^in[16]^in[20]^in[23]^in[24]^in[28]^in[30]^in[32]^in[37]^in[38]^in[39]^in[41]^in[48]^in[49]^in[52]^in[55]^in[56]^in[57]^in[60]^in[61]^in[62];//26 inputs
        syndrom[7] = in[ 2]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[13]^in[18]^in[19]^in[22]^in[25]^in[27]^in[31]^in[32]^in[37]^in[38]^in[42]^in[43]^in[46]^in[47]^in[51]^in[55]^in[56]^in[58]^in[59]^in[62]^in[63];//26 inputs
        extended_hamming_code_72_64_f = syndrom;
    end
endfunction
wire [8-1:0] stored_data_edc = extended_hamming_code_72_64_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_64_min_width (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [64-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_72_64_f
//Compute 8 bits Error Detection Code from a 64 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[0]: x   xx    xx   xx   x x  x  xx    xx  x x  x   x  xx  x x  xxxx  (26 inputs)
//  syndrom[1]: x   x x  x  xx   x  xx    xx   xx   x  xx    x xx    xx x x xxx  (26 inputs)
//  syndrom[2]: x    xx x    xx x    xx x    xx  x  xx    x x x   x xx   xxx x x (26 inputs)
//  syndrom[3]:  xx    x xx    x xx    x xx    x xx     xxx x     x xx   xxx  xx (26 inputs)
//  syndrom[4]:  x x   xx   x x  x x   xx   xx    xxx      xxx  xx    x  xxxx  x (26 inputs)
//  syndrom[5]:  x  xx    xx  x   xx x    xx  x  x x   x x   xx  x x   xxx  xx x (26 inputs)
//  syndrom[6]:   xx  x  x x   xx   x  xx   x x x    xxx x      xx  x  xxx  xxx  (26 inputs)
//  syndrom[7]:   xx   xx   xx    xx  x  x x   xx    xx   xx  xx   x   xx xx  xx (26 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 6 7)
//  input bit  3 used 3 times (syndrom bits 4 6 7)
//  input bit  4 used 3 times (syndrom bits 0 1 5)
//  input bit  5 used 3 times (syndrom bits 0 2 5)
//  input bit  6 used 3 times (syndrom bits 1 2 6)
//  input bit  7 used 3 times (syndrom bits 3 4 7)
//  input bit  8 used 3 times (syndrom bits 2 4 7)
//  input bit  9 used 3 times (syndrom bits 1 3 6)
//  input bit 10 used 3 times (syndrom bits 0 3 5)
//  input bit 11 used 3 times (syndrom bits 0 5 6)
//  input bit 12 used 3 times (syndrom bits 1 4 7)
//  input bit 13 used 3 times (syndrom bits 1 2 7)
//  input bit 14 used 3 times (syndrom bits 2 4 5)
//  input bit 15 used 3 times (syndrom bits 0 3 6)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 1 3 4)
//  input bit 18 used 3 times (syndrom bits 3 5 7)
//  input bit 19 used 3 times (syndrom bits 4 5 7)
//  input bit 20 used 3 times (syndrom bits 0 1 6)
//  input bit 21 used 3 times (syndrom bits 1 2 5)
//  input bit 22 used 3 times (syndrom bits 0 2 7)
//  input bit 23 used 3 times (syndrom bits 3 4 6)
//  input bit 24 used 3 times (syndrom bits 2 4 6)
//  input bit 25 used 3 times (syndrom bits 0 3 7)
//  input bit 26 used 3 times (syndrom bits 1 3 5)
//  input bit 27 used 3 times (syndrom bits 1 5 7)
//  input bit 28 used 3 times (syndrom bits 0 4 6)
//  input bit 29 used 3 times (syndrom bits 0 2 4)
//  input bit 30 used 3 times (syndrom bits 2 5 6)
//  input bit 31 used 3 times (syndrom bits 1 3 7)
//  input bit 32 used 3 times (syndrom bits 1 6 7)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 3 4)
//  input bit 35 used 3 times (syndrom bits 0 4 5)
//  input bit 36 used 3 times (syndrom bits 1 2 4)
//  input bit 37 used 3 times (syndrom bits 2 6 7)
//  input bit 38 used 3 times (syndrom bits 0 6 7)
//  input bit 39 used 3 times (syndrom bits 1 5 6)
//  input bit 40 used 3 times (syndrom bits 0 1 3)
//  input bit 41 used 3 times (syndrom bits 3 5 6)
//  input bit 42 used 3 times (syndrom bits 2 3 7)
//  input bit 43 used 3 times (syndrom bits 0 4 7)
//  input bit 44 used 3 times (syndrom bits 2 3 4)
//  input bit 45 used 3 times (syndrom bits 1 4 5)
//  input bit 46 used 3 times (syndrom bits 2 5 7)
//  input bit 47 used 3 times (syndrom bits 0 1 7)
//  input bit 48 used 3 times (syndrom bits 1 4 6)
//  input bit 49 used 3 times (syndrom bits 4 5 6)
//  input bit 50 used 3 times (syndrom bits 0 2 3)
//  input bit 51 used 3 times (syndrom bits 0 5 7)
//  input bit 52 used 3 times (syndrom bits 2 3 6)
//  input bit 53 used 3 times (syndrom bits 1 2 3)
//  input bit 54 used 3 times (syndrom bits 0 1 4)
//  input bit 55 used 3 times (syndrom bits 5 6 7)
//  input bit 56 used 5 times (syndrom bits 0 1 5 6 7)
//  input bit 57 used 5 times (syndrom bits 2 3 4 5 6)
//  input bit 58 used 5 times (syndrom bits 1 2 3 4 7)
//  input bit 59 used 5 times (syndrom bits 0 2 3 4 7)
//  input bit 60 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 61 used 5 times (syndrom bits 0 1 2 5 6)
//  input bit 62 used 5 times (syndrom bits 0 1 3 6 7)
//  input bit 63 used 5 times (syndrom bits 2 3 4 5 7)
function [8-1:0] extended_hamming_code_72_64_f;
    input [64-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 5]^in[10]^in[11]^in[15]^in[16]^in[20]^in[22]^in[25]^in[28]^in[29]^in[34]^in[35]^in[38]^in[40]^in[43]^in[47]^in[50]^in[51]^in[54]^in[56]^in[59]^in[60]^in[61]^in[62];//26 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 6]^in[ 9]^in[12]^in[13]^in[17]^in[20]^in[21]^in[26]^in[27]^in[31]^in[32]^in[36]^in[39]^in[40]^in[45]^in[47]^in[48]^in[53]^in[54]^in[56]^in[58]^in[60]^in[61]^in[62];//26 inputs
        syndrom[2] = in[ 0]^in[ 5]^in[ 6]^in[ 8]^in[13]^in[14]^in[16]^in[21]^in[22]^in[24]^in[29]^in[30]^in[33]^in[36]^in[37]^in[42]^in[44]^in[46]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[61]^in[63];//26 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 7]^in[ 9]^in[10]^in[15]^in[17]^in[18]^in[23]^in[25]^in[26]^in[31]^in[33]^in[34]^in[40]^in[41]^in[42]^in[44]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[62]^in[63];//26 inputs
        syndrom[4] = in[ 1]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[14]^in[17]^in[19]^in[23]^in[24]^in[28]^in[29]^in[34]^in[35]^in[36]^in[43]^in[44]^in[45]^in[48]^in[49]^in[54]^in[57]^in[58]^in[59]^in[60]^in[63];//26 inputs
        syndrom[5] = in[ 1]^in[ 4]^in[ 5]^in[10]^in[11]^in[14]^in[18]^in[19]^in[21]^in[26]^in[27]^in[30]^in[33]^in[35]^in[39]^in[41]^in[45]^in[46]^in[49]^in[51]^in[55]^in[56]^in[57]^in[60]^in[61]^in[63];//26 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 6]^in[ 9]^in[11]^in[15]^in[16]^in[20]^in[23]^in[24]^in[28]^in[30]^in[32]^in[37]^in[38]^in[39]^in[41]^in[48]^in[49]^in[52]^in[55]^in[56]^in[57]^in[60]^in[61]^in[62];//26 inputs
        syndrom[7] = in[ 2]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[13]^in[18]^in[19]^in[22]^in[25]^in[27]^in[31]^in[32]^in[37]^in[38]^in[42]^in[43]^in[46]^in[47]^in[51]^in[55]^in[56]^in[58]^in[59]^in[62]^in[63];//26 inputs
        extended_hamming_code_72_64_f = syndrom;
    end
endfunction
function [2+64-1:0] extended_hamming_code_72_64_f_correction_pattern_f;
    input [8-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [64-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {64{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			8'b00000000: begin
				correctable_error = 1'b0;
				correction_pattern = {64{1'b0}};
			end	
			8'b00000111: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 0]=1'b1;
			end
			8'b00111000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 1]=1'b1;
			end
			8'b11001000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 2]=1'b1;
			end
			8'b11010000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 3]=1'b1;
			end
			8'b00100011: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 4]=1'b1;
			end
			8'b00100101: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 5]=1'b1;
			end
			8'b01000110: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 6]=1'b1;
			end
			8'b10011000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 7]=1'b1;
			end
			8'b10010100: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 8]=1'b1;
			end
			8'b01001010: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 9]=1'b1;
			end
			8'b00101001: begin
				correction_pattern = {64{1'b0}};correction_pattern[10]=1'b1;
			end
			8'b01100001: begin
				correction_pattern = {64{1'b0}};correction_pattern[11]=1'b1;
			end
			8'b10010010: begin
				correction_pattern = {64{1'b0}};correction_pattern[12]=1'b1;
			end
			8'b10000110: begin
				correction_pattern = {64{1'b0}};correction_pattern[13]=1'b1;
			end
			8'b00110100: begin
				correction_pattern = {64{1'b0}};correction_pattern[14]=1'b1;
			end
			8'b01001001: begin
				correction_pattern = {64{1'b0}};correction_pattern[15]=1'b1;
			end
			8'b01000101: begin
				correction_pattern = {64{1'b0}};correction_pattern[16]=1'b1;
			end
			8'b00011010: begin
				correction_pattern = {64{1'b0}};correction_pattern[17]=1'b1;
			end
			8'b10101000: begin
				correction_pattern = {64{1'b0}};correction_pattern[18]=1'b1;
			end
			8'b10110000: begin
				correction_pattern = {64{1'b0}};correction_pattern[19]=1'b1;
			end
			8'b01000011: begin
				correction_pattern = {64{1'b0}};correction_pattern[20]=1'b1;
			end
			8'b00100110: begin
				correction_pattern = {64{1'b0}};correction_pattern[21]=1'b1;
			end
			8'b10000101: begin
				correction_pattern = {64{1'b0}};correction_pattern[22]=1'b1;
			end
			8'b01011000: begin
				correction_pattern = {64{1'b0}};correction_pattern[23]=1'b1;
			end
			8'b01010100: begin
				correction_pattern = {64{1'b0}};correction_pattern[24]=1'b1;
			end
			8'b10001001: begin
				correction_pattern = {64{1'b0}};correction_pattern[25]=1'b1;
			end
			8'b00101010: begin
				correction_pattern = {64{1'b0}};correction_pattern[26]=1'b1;
			end
			8'b10100010: begin
				correction_pattern = {64{1'b0}};correction_pattern[27]=1'b1;
			end
			8'b01010001: begin
				correction_pattern = {64{1'b0}};correction_pattern[28]=1'b1;
			end
			8'b00010101: begin
				correction_pattern = {64{1'b0}};correction_pattern[29]=1'b1;
			end
			8'b01100100: begin
				correction_pattern = {64{1'b0}};correction_pattern[30]=1'b1;
			end
			8'b10001010: begin
				correction_pattern = {64{1'b0}};correction_pattern[31]=1'b1;
			end
			8'b11000010: begin
				correction_pattern = {64{1'b0}};correction_pattern[32]=1'b1;
			end
			8'b00101100: begin
				correction_pattern = {64{1'b0}};correction_pattern[33]=1'b1;
			end
			8'b00011001: begin
				correction_pattern = {64{1'b0}};correction_pattern[34]=1'b1;
			end
			8'b00110001: begin
				correction_pattern = {64{1'b0}};correction_pattern[35]=1'b1;
			end
			8'b00010110: begin
				correction_pattern = {64{1'b0}};correction_pattern[36]=1'b1;
			end
			8'b11000100: begin
				correction_pattern = {64{1'b0}};correction_pattern[37]=1'b1;
			end
			8'b11000001: begin
				correction_pattern = {64{1'b0}};correction_pattern[38]=1'b1;
			end
			8'b01100010: begin
				correction_pattern = {64{1'b0}};correction_pattern[39]=1'b1;
			end
			8'b00001011: begin
				correction_pattern = {64{1'b0}};correction_pattern[40]=1'b1;
			end
			8'b01101000: begin
				correction_pattern = {64{1'b0}};correction_pattern[41]=1'b1;
			end
			8'b10001100: begin
				correction_pattern = {64{1'b0}};correction_pattern[42]=1'b1;
			end
			8'b10010001: begin
				correction_pattern = {64{1'b0}};correction_pattern[43]=1'b1;
			end
			8'b00011100: begin
				correction_pattern = {64{1'b0}};correction_pattern[44]=1'b1;
			end
			8'b00110010: begin
				correction_pattern = {64{1'b0}};correction_pattern[45]=1'b1;
			end
			8'b10100100: begin
				correction_pattern = {64{1'b0}};correction_pattern[46]=1'b1;
			end
			8'b10000011: begin
				correction_pattern = {64{1'b0}};correction_pattern[47]=1'b1;
			end
			8'b01010010: begin
				correction_pattern = {64{1'b0}};correction_pattern[48]=1'b1;
			end
			8'b01110000: begin
				correction_pattern = {64{1'b0}};correction_pattern[49]=1'b1;
			end
			8'b00001101: begin
				correction_pattern = {64{1'b0}};correction_pattern[50]=1'b1;
			end
			8'b10100001: begin
				correction_pattern = {64{1'b0}};correction_pattern[51]=1'b1;
			end
			8'b01001100: begin
				correction_pattern = {64{1'b0}};correction_pattern[52]=1'b1;
			end
			8'b00001110: begin
				correction_pattern = {64{1'b0}};correction_pattern[53]=1'b1;
			end
			8'b00010011: begin
				correction_pattern = {64{1'b0}};correction_pattern[54]=1'b1;
			end
			8'b11100000: begin
				correction_pattern = {64{1'b0}};correction_pattern[55]=1'b1;
			end
			8'b11100011: begin
				correction_pattern = {64{1'b0}};correction_pattern[56]=1'b1;
			end
			8'b01111100: begin
				correction_pattern = {64{1'b0}};correction_pattern[57]=1'b1;
			end
			8'b10011110: begin
				correction_pattern = {64{1'b0}};correction_pattern[58]=1'b1;
			end
			8'b10011101: begin
				correction_pattern = {64{1'b0}};correction_pattern[59]=1'b1;
			end
			8'b01110011: begin
				correction_pattern = {64{1'b0}};correction_pattern[60]=1'b1;
			end
			8'b01100111: begin
				correction_pattern = {64{1'b0}};correction_pattern[61]=1'b1;
			end
			8'b11001011: begin
				correction_pattern = {64{1'b0}};correction_pattern[62]=1'b1;
			end
			8'b10111100: begin
				correction_pattern = {64{1'b0}};correction_pattern[63]=1'b1;
			end
			8'b00000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b01000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b10000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_72_64_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [8-1:0] stored_data_edc = extended_hamming_code_72_64_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [64-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_72_64_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_96_min_width (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [7-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [7-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_103_96_f
//Compute 7 bits Error Detection Code from a 96 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 4 6)
//  input bit  4 used 2 times (syndrom bits 5 6)
//  input bit  5 used 2 times (syndrom bits 0 2)
//  input bit  6 used 2 times (syndrom bits 1 3)
//  input bit  7 used 2 times (syndrom bits 0 3)
//  input bit  8 used 2 times (syndrom bits 1 2)
//  input bit  9 used 2 times (syndrom bits 1 6)
//  input bit 10 used 2 times (syndrom bits 2 5)
//  input bit 11 used 2 times (syndrom bits 3 4)
//  input bit 12 used 2 times (syndrom bits 0 4)
//  input bit 13 used 2 times (syndrom bits 0 5)
//  input bit 14 used 2 times (syndrom bits 3 6)
//  input bit 15 used 2 times (syndrom bits 2 6)
//  input bit 16 used 2 times (syndrom bits 1 5)
//  input bit 17 used 2 times (syndrom bits 1 4)
//  input bit 18 used 2 times (syndrom bits 2 4)
//  input bit 19 used 2 times (syndrom bits 3 5)
//  input bit 20 used 2 times (syndrom bits 0 6)
//  input bit 21 used 3 times (syndrom bits 0 5 6)
//  input bit 22 used 3 times (syndrom bits 2 3 4)
//  input bit 23 used 3 times (syndrom bits 1 3 4)
//  input bit 24 used 3 times (syndrom bits 1 2 6)
//  input bit 25 used 3 times (syndrom bits 0 1 5)
//  input bit 26 used 3 times (syndrom bits 0 2 5)
//  input bit 27 used 3 times (syndrom bits 3 4 6)
//  input bit 28 used 3 times (syndrom bits 0 3 6)
//  input bit 29 used 3 times (syndrom bits 2 4 5)
//  input bit 30 used 3 times (syndrom bits 1 4 5)
//  input bit 31 used 3 times (syndrom bits 1 2 3)
//  input bit 32 used 3 times (syndrom bits 0 1 6)
//  input bit 33 used 3 times (syndrom bits 0 2 6)
//  input bit 34 used 3 times (syndrom bits 3 4 5)
//  input bit 35 used 3 times (syndrom bits 0 3 4)
//  input bit 36 used 3 times (syndrom bits 2 5 6)
//  input bit 37 used 3 times (syndrom bits 1 5 6)
//  input bit 38 used 3 times (syndrom bits 1 2 4)
//  input bit 39 used 3 times (syndrom bits 0 1 3)
//  input bit 40 used 3 times (syndrom bits 0 2 3)
//  input bit 41 used 3 times (syndrom bits 4 5 6)
//  input bit 42 used 3 times (syndrom bits 0 4 5)
//  input bit 43 used 3 times (syndrom bits 2 3 6)
//  input bit 44 used 3 times (syndrom bits 1 3 6)
//  input bit 45 used 3 times (syndrom bits 1 2 5)
//  input bit 46 used 3 times (syndrom bits 0 1 4)
//  input bit 47 used 3 times (syndrom bits 0 2 4)
//  input bit 48 used 3 times (syndrom bits 3 5 6)
//  input bit 49 used 3 times (syndrom bits 0 3 5)
//  input bit 50 used 3 times (syndrom bits 2 4 6)
//  input bit 51 used 3 times (syndrom bits 1 4 6)
//  input bit 52 used 3 times (syndrom bits 0 1 2)
//  input bit 53 used 3 times (syndrom bits 1 3 5)
//  input bit 54 used 3 times (syndrom bits 2 3 5)
//  input bit 55 used 3 times (syndrom bits 0 4 6)
//  input bit 56 used 4 times (syndrom bits 0 4 5 6)
//  input bit 57 used 4 times (syndrom bits 0 1 2 3)
//  input bit 58 used 4 times (syndrom bits 1 2 3 6)
//  input bit 59 used 4 times (syndrom bits 2 3 4 5)
//  input bit 60 used 4 times (syndrom bits 1 4 5 6)
//  input bit 61 used 4 times (syndrom bits 0 1 4 5)
//  input bit 62 used 4 times (syndrom bits 0 2 3 6)
//  input bit 63 used 4 times (syndrom bits 0 3 4 6)
//  input bit 64 used 4 times (syndrom bits 0 1 2 5)
//  input bit 65 used 4 times (syndrom bits 1 2 5 6)
//  input bit 66 used 4 times (syndrom bits 1 2 3 4)
//  input bit 67 used 4 times (syndrom bits 3 4 5 6)
//  input bit 68 used 4 times (syndrom bits 0 3 4 5)
//  input bit 69 used 4 times (syndrom bits 0 1 2 6)
//  input bit 70 used 4 times (syndrom bits 0 2 4 6)
//  input bit 71 used 4 times (syndrom bits 0 1 3 5)
//  input bit 72 used 4 times (syndrom bits 1 3 5 6)
//  input bit 73 used 4 times (syndrom bits 1 2 4 5)
//  input bit 74 used 4 times (syndrom bits 2 3 4 6)
//  input bit 75 used 4 times (syndrom bits 0 2 3 4)
//  input bit 76 used 4 times (syndrom bits 0 1 5 6)
//  input bit 77 used 4 times (syndrom bits 0 1 4 6)
//  input bit 78 used 4 times (syndrom bits 0 2 3 5)
//  input bit 79 used 4 times (syndrom bits 2 3 5 6)
//  input bit 80 used 4 times (syndrom bits 1 3 4 5)
//  input bit 81 used 4 times (syndrom bits 1 2 4 6)
//  input bit 82 used 4 times (syndrom bits 0 1 2 4)
//  input bit 83 used 4 times (syndrom bits 0 3 5 6)
//  input bit 84 used 4 times (syndrom bits 0 2 5 6)
//  input bit 85 used 4 times (syndrom bits 0 1 3 4)
//  input bit 86 used 4 times (syndrom bits 1 3 4 6)
//  input bit 87 used 4 times (syndrom bits 1 2 3 5)
//  input bit 88 used 4 times (syndrom bits 2 4 5 6)
//  input bit 89 used 4 times (syndrom bits 0 2 4 5)
//  input bit 90 used 4 times (syndrom bits 0 1 3 6)
//  input bit 91 used 5 times (syndrom bits 0 1 3 5 6)
//  input bit 92 used 5 times (syndrom bits 0 2 3 4 6)
//  input bit 93 used 5 times (syndrom bits 0 1 2 4 5)
//  input bit 94 used 5 times (syndrom bits 1 2 4 5 6)
//  input bit 95 used 5 times (syndrom bits 1 2 3 4 5)
function [7-1:0] hamming_code_103_96_f;
    input [96-1:0] in;
    reg [7-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 5]^in[ 7]^in[12]^in[13]^in[20]^in[21]^in[25]^in[26]^in[28]^in[32]^in[33]^in[35]^in[39]^in[40]^in[42]^in[46]^in[47]^in[49]^in[52]^in[55]^in[56]^in[57]^in[61]^in[62]^in[63]^in[64]^in[68]^in[69]^in[70]^in[71]^in[75]^in[76]^in[77]^in[78]^in[82]^in[83]^in[84]^in[85]^in[89]^in[90]^in[91]^in[92]^in[93];//44 inputs
        syndrom[1] = in[ 0]^in[ 6]^in[ 8]^in[ 9]^in[16]^in[17]^in[23]^in[24]^in[25]^in[30]^in[31]^in[32]^in[37]^in[38]^in[39]^in[44]^in[45]^in[46]^in[51]^in[52]^in[53]^in[57]^in[58]^in[60]^in[61]^in[64]^in[65]^in[66]^in[69]^in[71]^in[72]^in[73]^in[76]^in[77]^in[80]^in[81]^in[82]^in[85]^in[86]^in[87]^in[90]^in[91]^in[93]^in[94]^in[95];//45 inputs
        syndrom[2] = in[ 1]^in[ 5]^in[ 8]^in[10]^in[15]^in[18]^in[22]^in[24]^in[26]^in[29]^in[31]^in[33]^in[36]^in[38]^in[40]^in[43]^in[45]^in[47]^in[50]^in[52]^in[54]^in[57]^in[58]^in[59]^in[62]^in[64]^in[65]^in[66]^in[69]^in[70]^in[73]^in[74]^in[75]^in[78]^in[79]^in[81]^in[82]^in[84]^in[87]^in[88]^in[89]^in[92]^in[93]^in[94]^in[95];//45 inputs
        syndrom[3] = in[ 1]^in[ 6]^in[ 7]^in[11]^in[14]^in[19]^in[22]^in[23]^in[27]^in[28]^in[31]^in[34]^in[35]^in[39]^in[40]^in[43]^in[44]^in[48]^in[49]^in[53]^in[54]^in[57]^in[58]^in[59]^in[62]^in[63]^in[66]^in[67]^in[68]^in[71]^in[72]^in[74]^in[75]^in[78]^in[79]^in[80]^in[83]^in[85]^in[86]^in[87]^in[90]^in[91]^in[92]^in[95];//44 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[11]^in[12]^in[17]^in[18]^in[22]^in[23]^in[27]^in[29]^in[30]^in[34]^in[35]^in[38]^in[41]^in[42]^in[46]^in[47]^in[50]^in[51]^in[55]^in[56]^in[59]^in[60]^in[61]^in[63]^in[66]^in[67]^in[68]^in[70]^in[73]^in[74]^in[75]^in[77]^in[80]^in[81]^in[82]^in[85]^in[86]^in[88]^in[89]^in[92]^in[93]^in[94]^in[95];//45 inputs
        syndrom[5] = in[ 2]^in[ 4]^in[10]^in[13]^in[16]^in[19]^in[21]^in[25]^in[26]^in[29]^in[30]^in[34]^in[36]^in[37]^in[41]^in[42]^in[45]^in[48]^in[49]^in[53]^in[54]^in[56]^in[59]^in[60]^in[61]^in[64]^in[65]^in[67]^in[68]^in[71]^in[72]^in[73]^in[76]^in[78]^in[79]^in[80]^in[83]^in[84]^in[87]^in[88]^in[89]^in[91]^in[93]^in[94]^in[95];//45 inputs
        syndrom[6] = in[ 3]^in[ 4]^in[ 9]^in[14]^in[15]^in[20]^in[21]^in[24]^in[27]^in[28]^in[32]^in[33]^in[36]^in[37]^in[41]^in[43]^in[44]^in[48]^in[50]^in[51]^in[55]^in[56]^in[58]^in[60]^in[62]^in[63]^in[65]^in[67]^in[69]^in[70]^in[72]^in[74]^in[76]^in[77]^in[79]^in[81]^in[83]^in[84]^in[86]^in[88]^in[90]^in[91]^in[92]^in[94];//44 inputs
        hamming_code_103_96_f = syndrom;
    end
endfunction
wire [7-1:0] stored_data_edc = hamming_code_103_96_f(i_stored_data);
wire [7-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_96_min_width (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_104_96_f
//Compute 8 bits Error Detection Code from a 96 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 6 7)
//  input bit  3 used 3 times (syndrom bits 4 6 7)
//  input bit  4 used 3 times (syndrom bits 0 1 5)
//  input bit  5 used 3 times (syndrom bits 0 2 5)
//  input bit  6 used 3 times (syndrom bits 1 2 6)
//  input bit  7 used 3 times (syndrom bits 3 4 7)
//  input bit  8 used 3 times (syndrom bits 2 4 7)
//  input bit  9 used 3 times (syndrom bits 1 3 6)
//  input bit 10 used 3 times (syndrom bits 0 3 5)
//  input bit 11 used 3 times (syndrom bits 0 5 6)
//  input bit 12 used 3 times (syndrom bits 1 4 7)
//  input bit 13 used 3 times (syndrom bits 1 2 7)
//  input bit 14 used 3 times (syndrom bits 2 4 5)
//  input bit 15 used 3 times (syndrom bits 0 3 6)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 1 3 4)
//  input bit 18 used 3 times (syndrom bits 3 5 7)
//  input bit 19 used 3 times (syndrom bits 4 5 7)
//  input bit 20 used 3 times (syndrom bits 0 1 6)
//  input bit 21 used 3 times (syndrom bits 1 2 5)
//  input bit 22 used 3 times (syndrom bits 0 2 7)
//  input bit 23 used 3 times (syndrom bits 3 4 6)
//  input bit 24 used 3 times (syndrom bits 2 4 6)
//  input bit 25 used 3 times (syndrom bits 0 3 7)
//  input bit 26 used 3 times (syndrom bits 1 3 5)
//  input bit 27 used 3 times (syndrom bits 1 5 7)
//  input bit 28 used 3 times (syndrom bits 0 4 6)
//  input bit 29 used 3 times (syndrom bits 0 2 4)
//  input bit 30 used 3 times (syndrom bits 2 5 6)
//  input bit 31 used 3 times (syndrom bits 1 3 7)
//  input bit 32 used 3 times (syndrom bits 1 6 7)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 3 4)
//  input bit 35 used 3 times (syndrom bits 0 4 5)
//  input bit 36 used 3 times (syndrom bits 1 2 4)
//  input bit 37 used 3 times (syndrom bits 2 6 7)
//  input bit 38 used 3 times (syndrom bits 0 6 7)
//  input bit 39 used 3 times (syndrom bits 1 5 6)
//  input bit 40 used 3 times (syndrom bits 0 1 3)
//  input bit 41 used 3 times (syndrom bits 3 5 6)
//  input bit 42 used 3 times (syndrom bits 2 3 7)
//  input bit 43 used 3 times (syndrom bits 0 4 7)
//  input bit 44 used 3 times (syndrom bits 2 3 4)
//  input bit 45 used 3 times (syndrom bits 1 4 5)
//  input bit 46 used 3 times (syndrom bits 2 5 7)
//  input bit 47 used 3 times (syndrom bits 0 1 7)
//  input bit 48 used 3 times (syndrom bits 1 4 6)
//  input bit 49 used 3 times (syndrom bits 4 5 6)
//  input bit 50 used 3 times (syndrom bits 0 2 3)
//  input bit 51 used 3 times (syndrom bits 0 5 7)
//  input bit 52 used 3 times (syndrom bits 2 3 6)
//  input bit 53 used 3 times (syndrom bits 1 2 3)
//  input bit 54 used 3 times (syndrom bits 0 1 4)
//  input bit 55 used 3 times (syndrom bits 5 6 7)
//  input bit 56 used 5 times (syndrom bits 0 1 5 6 7)
//  input bit 57 used 5 times (syndrom bits 2 3 4 5 6)
//  input bit 58 used 5 times (syndrom bits 1 2 3 4 7)
//  input bit 59 used 5 times (syndrom bits 0 2 3 4 7)
//  input bit 60 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 61 used 5 times (syndrom bits 0 1 2 5 6)
//  input bit 62 used 5 times (syndrom bits 0 1 3 6 7)
//  input bit 63 used 5 times (syndrom bits 2 3 4 5 7)
//  input bit 64 used 5 times (syndrom bits 0 2 3 5 7)
//  input bit 65 used 5 times (syndrom bits 1 3 4 6 7)
//  input bit 66 used 5 times (syndrom bits 1 2 4 5 6)
//  input bit 67 used 5 times (syndrom bits 0 1 2 4 6)
//  input bit 68 used 5 times (syndrom bits 0 3 4 5 7)
//  input bit 69 used 5 times (syndrom bits 0 1 3 5 7)
//  input bit 70 used 5 times (syndrom bits 0 2 3 5 6)
//  input bit 71 used 5 times (syndrom bits 1 2 4 6 7)
//  input bit 72 used 5 times (syndrom bits 0 1 2 6 7)
//  input bit 73 used 5 times (syndrom bits 3 4 5 6 7)
//  input bit 74 used 5 times (syndrom bits 1 2 3 4 5)
//  input bit 75 used 5 times (syndrom bits 0 2 3 4 5)
//  input bit 76 used 5 times (syndrom bits 0 1 4 6 7)
//  input bit 77 used 5 times (syndrom bits 0 1 3 5 6)
//  input bit 78 used 5 times (syndrom bits 0 1 2 5 7)
//  input bit 79 used 5 times (syndrom bits 2 3 4 6 7)
//  input bit 80 used 5 times (syndrom bits 0 2 3 6 7)
//  input bit 81 used 5 times (syndrom bits 1 2 4 5 7)
//  input bit 82 used 5 times (syndrom bits 1 3 4 5 6)
//  input bit 83 used 5 times (syndrom bits 0 1 3 4 5)
//  input bit 84 used 5 times (syndrom bits 0 2 4 6 7)
//  input bit 85 used 5 times (syndrom bits 0 2 5 6 7)
//  input bit 86 used 5 times (syndrom bits 0 1 2 3 6)
//  input bit 87 used 5 times (syndrom bits 1 3 4 5 7)
//  input bit 88 used 5 times (syndrom bits 1 3 5 6 7)
//  input bit 89 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 90 used 5 times (syndrom bits 0 2 4 5 7)
//  input bit 91 used 5 times (syndrom bits 0 2 4 5 6)
//  input bit 92 used 5 times (syndrom bits 1 2 3 6 7)
//  input bit 93 used 5 times (syndrom bits 1 4 5 6 7)
//  input bit 94 used 5 times (syndrom bits 0 3 4 6 7)
//  input bit 95 used 5 times (syndrom bits 0 1 2 3 5)
function [8-1:0] extended_hamming_code_104_96_f;
    input [96-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 5]^in[10]^in[11]^in[15]^in[16]^in[20]^in[22]^in[25]^in[28]^in[29]^in[34]^in[35]^in[38]^in[40]^in[43]^in[47]^in[50]^in[51]^in[54]^in[56]^in[59]^in[60]^in[61]^in[62]^in[64]^in[67]^in[68]^in[69]^in[70]^in[72]^in[75]^in[76]^in[77]^in[78]^in[80]^in[83]^in[84]^in[85]^in[86]^in[89]^in[90]^in[91]^in[94]^in[95];//46 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 6]^in[ 9]^in[12]^in[13]^in[17]^in[20]^in[21]^in[26]^in[27]^in[31]^in[32]^in[36]^in[39]^in[40]^in[45]^in[47]^in[48]^in[53]^in[54]^in[56]^in[58]^in[60]^in[61]^in[62]^in[65]^in[66]^in[67]^in[69]^in[71]^in[72]^in[74]^in[76]^in[77]^in[78]^in[81]^in[82]^in[83]^in[86]^in[87]^in[88]^in[89]^in[92]^in[93]^in[95];//46 inputs
        syndrom[2] = in[ 0]^in[ 5]^in[ 6]^in[ 8]^in[13]^in[14]^in[16]^in[21]^in[22]^in[24]^in[29]^in[30]^in[33]^in[36]^in[37]^in[42]^in[44]^in[46]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[61]^in[63]^in[64]^in[66]^in[67]^in[70]^in[71]^in[72]^in[74]^in[75]^in[78]^in[79]^in[80]^in[81]^in[84]^in[85]^in[86]^in[89]^in[90]^in[91]^in[92]^in[95];//46 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 7]^in[ 9]^in[10]^in[15]^in[17]^in[18]^in[23]^in[25]^in[26]^in[31]^in[33]^in[34]^in[40]^in[41]^in[42]^in[44]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[62]^in[63]^in[64]^in[65]^in[68]^in[69]^in[70]^in[73]^in[74]^in[75]^in[77]^in[79]^in[80]^in[82]^in[83]^in[86]^in[87]^in[88]^in[89]^in[92]^in[94]^in[95];//46 inputs
        syndrom[4] = in[ 1]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[14]^in[17]^in[19]^in[23]^in[24]^in[28]^in[29]^in[34]^in[35]^in[36]^in[43]^in[44]^in[45]^in[48]^in[49]^in[54]^in[57]^in[58]^in[59]^in[60]^in[63]^in[65]^in[66]^in[67]^in[68]^in[71]^in[73]^in[74]^in[75]^in[76]^in[79]^in[81]^in[82]^in[83]^in[84]^in[87]^in[89]^in[90]^in[91]^in[93]^in[94];//46 inputs
        syndrom[5] = in[ 1]^in[ 4]^in[ 5]^in[10]^in[11]^in[14]^in[18]^in[19]^in[21]^in[26]^in[27]^in[30]^in[33]^in[35]^in[39]^in[41]^in[45]^in[46]^in[49]^in[51]^in[55]^in[56]^in[57]^in[60]^in[61]^in[63]^in[64]^in[66]^in[68]^in[69]^in[70]^in[73]^in[74]^in[75]^in[77]^in[78]^in[81]^in[82]^in[83]^in[85]^in[87]^in[88]^in[90]^in[91]^in[93]^in[95];//46 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 6]^in[ 9]^in[11]^in[15]^in[16]^in[20]^in[23]^in[24]^in[28]^in[30]^in[32]^in[37]^in[38]^in[39]^in[41]^in[48]^in[49]^in[52]^in[55]^in[56]^in[57]^in[60]^in[61]^in[62]^in[65]^in[66]^in[67]^in[70]^in[71]^in[72]^in[73]^in[76]^in[77]^in[79]^in[80]^in[82]^in[84]^in[85]^in[86]^in[88]^in[91]^in[92]^in[93]^in[94];//46 inputs
        syndrom[7] = in[ 2]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[13]^in[18]^in[19]^in[22]^in[25]^in[27]^in[31]^in[32]^in[37]^in[38]^in[42]^in[43]^in[46]^in[47]^in[51]^in[55]^in[56]^in[58]^in[59]^in[62]^in[63]^in[64]^in[65]^in[68]^in[69]^in[71]^in[72]^in[73]^in[76]^in[78]^in[79]^in[80]^in[81]^in[84]^in[85]^in[87]^in[88]^in[90]^in[92]^in[93]^in[94];//46 inputs
        extended_hamming_code_104_96_f = syndrom;
    end
endfunction
wire [8-1:0] stored_data_edc = extended_hamming_code_104_96_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_96_min_width (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [96-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_104_96_f
//Compute 8 bits Error Detection Code from a 96 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 6 7)
//  input bit  3 used 3 times (syndrom bits 4 6 7)
//  input bit  4 used 3 times (syndrom bits 0 1 5)
//  input bit  5 used 3 times (syndrom bits 0 2 5)
//  input bit  6 used 3 times (syndrom bits 1 2 6)
//  input bit  7 used 3 times (syndrom bits 3 4 7)
//  input bit  8 used 3 times (syndrom bits 2 4 7)
//  input bit  9 used 3 times (syndrom bits 1 3 6)
//  input bit 10 used 3 times (syndrom bits 0 3 5)
//  input bit 11 used 3 times (syndrom bits 0 5 6)
//  input bit 12 used 3 times (syndrom bits 1 4 7)
//  input bit 13 used 3 times (syndrom bits 1 2 7)
//  input bit 14 used 3 times (syndrom bits 2 4 5)
//  input bit 15 used 3 times (syndrom bits 0 3 6)
//  input bit 16 used 3 times (syndrom bits 0 2 6)
//  input bit 17 used 3 times (syndrom bits 1 3 4)
//  input bit 18 used 3 times (syndrom bits 3 5 7)
//  input bit 19 used 3 times (syndrom bits 4 5 7)
//  input bit 20 used 3 times (syndrom bits 0 1 6)
//  input bit 21 used 3 times (syndrom bits 1 2 5)
//  input bit 22 used 3 times (syndrom bits 0 2 7)
//  input bit 23 used 3 times (syndrom bits 3 4 6)
//  input bit 24 used 3 times (syndrom bits 2 4 6)
//  input bit 25 used 3 times (syndrom bits 0 3 7)
//  input bit 26 used 3 times (syndrom bits 1 3 5)
//  input bit 27 used 3 times (syndrom bits 1 5 7)
//  input bit 28 used 3 times (syndrom bits 0 4 6)
//  input bit 29 used 3 times (syndrom bits 0 2 4)
//  input bit 30 used 3 times (syndrom bits 2 5 6)
//  input bit 31 used 3 times (syndrom bits 1 3 7)
//  input bit 32 used 3 times (syndrom bits 1 6 7)
//  input bit 33 used 3 times (syndrom bits 2 3 5)
//  input bit 34 used 3 times (syndrom bits 0 3 4)
//  input bit 35 used 3 times (syndrom bits 0 4 5)
//  input bit 36 used 3 times (syndrom bits 1 2 4)
//  input bit 37 used 3 times (syndrom bits 2 6 7)
//  input bit 38 used 3 times (syndrom bits 0 6 7)
//  input bit 39 used 3 times (syndrom bits 1 5 6)
//  input bit 40 used 3 times (syndrom bits 0 1 3)
//  input bit 41 used 3 times (syndrom bits 3 5 6)
//  input bit 42 used 3 times (syndrom bits 2 3 7)
//  input bit 43 used 3 times (syndrom bits 0 4 7)
//  input bit 44 used 3 times (syndrom bits 2 3 4)
//  input bit 45 used 3 times (syndrom bits 1 4 5)
//  input bit 46 used 3 times (syndrom bits 2 5 7)
//  input bit 47 used 3 times (syndrom bits 0 1 7)
//  input bit 48 used 3 times (syndrom bits 1 4 6)
//  input bit 49 used 3 times (syndrom bits 4 5 6)
//  input bit 50 used 3 times (syndrom bits 0 2 3)
//  input bit 51 used 3 times (syndrom bits 0 5 7)
//  input bit 52 used 3 times (syndrom bits 2 3 6)
//  input bit 53 used 3 times (syndrom bits 1 2 3)
//  input bit 54 used 3 times (syndrom bits 0 1 4)
//  input bit 55 used 3 times (syndrom bits 5 6 7)
//  input bit 56 used 5 times (syndrom bits 0 1 5 6 7)
//  input bit 57 used 5 times (syndrom bits 2 3 4 5 6)
//  input bit 58 used 5 times (syndrom bits 1 2 3 4 7)
//  input bit 59 used 5 times (syndrom bits 0 2 3 4 7)
//  input bit 60 used 5 times (syndrom bits 0 1 4 5 6)
//  input bit 61 used 5 times (syndrom bits 0 1 2 5 6)
//  input bit 62 used 5 times (syndrom bits 0 1 3 6 7)
//  input bit 63 used 5 times (syndrom bits 2 3 4 5 7)
//  input bit 64 used 5 times (syndrom bits 0 2 3 5 7)
//  input bit 65 used 5 times (syndrom bits 1 3 4 6 7)
//  input bit 66 used 5 times (syndrom bits 1 2 4 5 6)
//  input bit 67 used 5 times (syndrom bits 0 1 2 4 6)
//  input bit 68 used 5 times (syndrom bits 0 3 4 5 7)
//  input bit 69 used 5 times (syndrom bits 0 1 3 5 7)
//  input bit 70 used 5 times (syndrom bits 0 2 3 5 6)
//  input bit 71 used 5 times (syndrom bits 1 2 4 6 7)
//  input bit 72 used 5 times (syndrom bits 0 1 2 6 7)
//  input bit 73 used 5 times (syndrom bits 3 4 5 6 7)
//  input bit 74 used 5 times (syndrom bits 1 2 3 4 5)
//  input bit 75 used 5 times (syndrom bits 0 2 3 4 5)
//  input bit 76 used 5 times (syndrom bits 0 1 4 6 7)
//  input bit 77 used 5 times (syndrom bits 0 1 3 5 6)
//  input bit 78 used 5 times (syndrom bits 0 1 2 5 7)
//  input bit 79 used 5 times (syndrom bits 2 3 4 6 7)
//  input bit 80 used 5 times (syndrom bits 0 2 3 6 7)
//  input bit 81 used 5 times (syndrom bits 1 2 4 5 7)
//  input bit 82 used 5 times (syndrom bits 1 3 4 5 6)
//  input bit 83 used 5 times (syndrom bits 0 1 3 4 5)
//  input bit 84 used 5 times (syndrom bits 0 2 4 6 7)
//  input bit 85 used 5 times (syndrom bits 0 2 5 6 7)
//  input bit 86 used 5 times (syndrom bits 0 1 2 3 6)
//  input bit 87 used 5 times (syndrom bits 1 3 4 5 7)
//  input bit 88 used 5 times (syndrom bits 1 3 5 6 7)
//  input bit 89 used 5 times (syndrom bits 0 1 2 3 4)
//  input bit 90 used 5 times (syndrom bits 0 2 4 5 7)
//  input bit 91 used 5 times (syndrom bits 0 2 4 5 6)
//  input bit 92 used 5 times (syndrom bits 1 2 3 6 7)
//  input bit 93 used 5 times (syndrom bits 1 4 5 6 7)
//  input bit 94 used 5 times (syndrom bits 0 3 4 6 7)
//  input bit 95 used 5 times (syndrom bits 0 1 2 3 5)
function [8-1:0] extended_hamming_code_104_96_f;
    input [96-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 5]^in[10]^in[11]^in[15]^in[16]^in[20]^in[22]^in[25]^in[28]^in[29]^in[34]^in[35]^in[38]^in[40]^in[43]^in[47]^in[50]^in[51]^in[54]^in[56]^in[59]^in[60]^in[61]^in[62]^in[64]^in[67]^in[68]^in[69]^in[70]^in[72]^in[75]^in[76]^in[77]^in[78]^in[80]^in[83]^in[84]^in[85]^in[86]^in[89]^in[90]^in[91]^in[94]^in[95];//46 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 6]^in[ 9]^in[12]^in[13]^in[17]^in[20]^in[21]^in[26]^in[27]^in[31]^in[32]^in[36]^in[39]^in[40]^in[45]^in[47]^in[48]^in[53]^in[54]^in[56]^in[58]^in[60]^in[61]^in[62]^in[65]^in[66]^in[67]^in[69]^in[71]^in[72]^in[74]^in[76]^in[77]^in[78]^in[81]^in[82]^in[83]^in[86]^in[87]^in[88]^in[89]^in[92]^in[93]^in[95];//46 inputs
        syndrom[2] = in[ 0]^in[ 5]^in[ 6]^in[ 8]^in[13]^in[14]^in[16]^in[21]^in[22]^in[24]^in[29]^in[30]^in[33]^in[36]^in[37]^in[42]^in[44]^in[46]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[61]^in[63]^in[64]^in[66]^in[67]^in[70]^in[71]^in[72]^in[74]^in[75]^in[78]^in[79]^in[80]^in[81]^in[84]^in[85]^in[86]^in[89]^in[90]^in[91]^in[92]^in[95];//46 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 7]^in[ 9]^in[10]^in[15]^in[17]^in[18]^in[23]^in[25]^in[26]^in[31]^in[33]^in[34]^in[40]^in[41]^in[42]^in[44]^in[50]^in[52]^in[53]^in[57]^in[58]^in[59]^in[62]^in[63]^in[64]^in[65]^in[68]^in[69]^in[70]^in[73]^in[74]^in[75]^in[77]^in[79]^in[80]^in[82]^in[83]^in[86]^in[87]^in[88]^in[89]^in[92]^in[94]^in[95];//46 inputs
        syndrom[4] = in[ 1]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[14]^in[17]^in[19]^in[23]^in[24]^in[28]^in[29]^in[34]^in[35]^in[36]^in[43]^in[44]^in[45]^in[48]^in[49]^in[54]^in[57]^in[58]^in[59]^in[60]^in[63]^in[65]^in[66]^in[67]^in[68]^in[71]^in[73]^in[74]^in[75]^in[76]^in[79]^in[81]^in[82]^in[83]^in[84]^in[87]^in[89]^in[90]^in[91]^in[93]^in[94];//46 inputs
        syndrom[5] = in[ 1]^in[ 4]^in[ 5]^in[10]^in[11]^in[14]^in[18]^in[19]^in[21]^in[26]^in[27]^in[30]^in[33]^in[35]^in[39]^in[41]^in[45]^in[46]^in[49]^in[51]^in[55]^in[56]^in[57]^in[60]^in[61]^in[63]^in[64]^in[66]^in[68]^in[69]^in[70]^in[73]^in[74]^in[75]^in[77]^in[78]^in[81]^in[82]^in[83]^in[85]^in[87]^in[88]^in[90]^in[91]^in[93]^in[95];//46 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 6]^in[ 9]^in[11]^in[15]^in[16]^in[20]^in[23]^in[24]^in[28]^in[30]^in[32]^in[37]^in[38]^in[39]^in[41]^in[48]^in[49]^in[52]^in[55]^in[56]^in[57]^in[60]^in[61]^in[62]^in[65]^in[66]^in[67]^in[70]^in[71]^in[72]^in[73]^in[76]^in[77]^in[79]^in[80]^in[82]^in[84]^in[85]^in[86]^in[88]^in[91]^in[92]^in[93]^in[94];//46 inputs
        syndrom[7] = in[ 2]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[13]^in[18]^in[19]^in[22]^in[25]^in[27]^in[31]^in[32]^in[37]^in[38]^in[42]^in[43]^in[46]^in[47]^in[51]^in[55]^in[56]^in[58]^in[59]^in[62]^in[63]^in[64]^in[65]^in[68]^in[69]^in[71]^in[72]^in[73]^in[76]^in[78]^in[79]^in[80]^in[81]^in[84]^in[85]^in[87]^in[88]^in[90]^in[92]^in[93]^in[94];//46 inputs
        extended_hamming_code_104_96_f = syndrom;
    end
endfunction
function [2+96-1:0] extended_hamming_code_104_96_f_correction_pattern_f;
    input [8-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [96-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {96{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			8'b00000000: begin
				correctable_error = 1'b0;
				correction_pattern = {96{1'b0}};
			end	
			8'b00000111: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 0]=1'b1;
			end
			8'b00111000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 1]=1'b1;
			end
			8'b11001000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 2]=1'b1;
			end
			8'b11010000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 3]=1'b1;
			end
			8'b00100011: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 4]=1'b1;
			end
			8'b00100101: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 5]=1'b1;
			end
			8'b01000110: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 6]=1'b1;
			end
			8'b10011000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 7]=1'b1;
			end
			8'b10010100: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 8]=1'b1;
			end
			8'b01001010: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 9]=1'b1;
			end
			8'b00101001: begin
				correction_pattern = {96{1'b0}};correction_pattern[10]=1'b1;
			end
			8'b01100001: begin
				correction_pattern = {96{1'b0}};correction_pattern[11]=1'b1;
			end
			8'b10010010: begin
				correction_pattern = {96{1'b0}};correction_pattern[12]=1'b1;
			end
			8'b10000110: begin
				correction_pattern = {96{1'b0}};correction_pattern[13]=1'b1;
			end
			8'b00110100: begin
				correction_pattern = {96{1'b0}};correction_pattern[14]=1'b1;
			end
			8'b01001001: begin
				correction_pattern = {96{1'b0}};correction_pattern[15]=1'b1;
			end
			8'b01000101: begin
				correction_pattern = {96{1'b0}};correction_pattern[16]=1'b1;
			end
			8'b00011010: begin
				correction_pattern = {96{1'b0}};correction_pattern[17]=1'b1;
			end
			8'b10101000: begin
				correction_pattern = {96{1'b0}};correction_pattern[18]=1'b1;
			end
			8'b10110000: begin
				correction_pattern = {96{1'b0}};correction_pattern[19]=1'b1;
			end
			8'b01000011: begin
				correction_pattern = {96{1'b0}};correction_pattern[20]=1'b1;
			end
			8'b00100110: begin
				correction_pattern = {96{1'b0}};correction_pattern[21]=1'b1;
			end
			8'b10000101: begin
				correction_pattern = {96{1'b0}};correction_pattern[22]=1'b1;
			end
			8'b01011000: begin
				correction_pattern = {96{1'b0}};correction_pattern[23]=1'b1;
			end
			8'b01010100: begin
				correction_pattern = {96{1'b0}};correction_pattern[24]=1'b1;
			end
			8'b10001001: begin
				correction_pattern = {96{1'b0}};correction_pattern[25]=1'b1;
			end
			8'b00101010: begin
				correction_pattern = {96{1'b0}};correction_pattern[26]=1'b1;
			end
			8'b10100010: begin
				correction_pattern = {96{1'b0}};correction_pattern[27]=1'b1;
			end
			8'b01010001: begin
				correction_pattern = {96{1'b0}};correction_pattern[28]=1'b1;
			end
			8'b00010101: begin
				correction_pattern = {96{1'b0}};correction_pattern[29]=1'b1;
			end
			8'b01100100: begin
				correction_pattern = {96{1'b0}};correction_pattern[30]=1'b1;
			end
			8'b10001010: begin
				correction_pattern = {96{1'b0}};correction_pattern[31]=1'b1;
			end
			8'b11000010: begin
				correction_pattern = {96{1'b0}};correction_pattern[32]=1'b1;
			end
			8'b00101100: begin
				correction_pattern = {96{1'b0}};correction_pattern[33]=1'b1;
			end
			8'b00011001: begin
				correction_pattern = {96{1'b0}};correction_pattern[34]=1'b1;
			end
			8'b00110001: begin
				correction_pattern = {96{1'b0}};correction_pattern[35]=1'b1;
			end
			8'b00010110: begin
				correction_pattern = {96{1'b0}};correction_pattern[36]=1'b1;
			end
			8'b11000100: begin
				correction_pattern = {96{1'b0}};correction_pattern[37]=1'b1;
			end
			8'b11000001: begin
				correction_pattern = {96{1'b0}};correction_pattern[38]=1'b1;
			end
			8'b01100010: begin
				correction_pattern = {96{1'b0}};correction_pattern[39]=1'b1;
			end
			8'b00001011: begin
				correction_pattern = {96{1'b0}};correction_pattern[40]=1'b1;
			end
			8'b01101000: begin
				correction_pattern = {96{1'b0}};correction_pattern[41]=1'b1;
			end
			8'b10001100: begin
				correction_pattern = {96{1'b0}};correction_pattern[42]=1'b1;
			end
			8'b10010001: begin
				correction_pattern = {96{1'b0}};correction_pattern[43]=1'b1;
			end
			8'b00011100: begin
				correction_pattern = {96{1'b0}};correction_pattern[44]=1'b1;
			end
			8'b00110010: begin
				correction_pattern = {96{1'b0}};correction_pattern[45]=1'b1;
			end
			8'b10100100: begin
				correction_pattern = {96{1'b0}};correction_pattern[46]=1'b1;
			end
			8'b10000011: begin
				correction_pattern = {96{1'b0}};correction_pattern[47]=1'b1;
			end
			8'b01010010: begin
				correction_pattern = {96{1'b0}};correction_pattern[48]=1'b1;
			end
			8'b01110000: begin
				correction_pattern = {96{1'b0}};correction_pattern[49]=1'b1;
			end
			8'b00001101: begin
				correction_pattern = {96{1'b0}};correction_pattern[50]=1'b1;
			end
			8'b10100001: begin
				correction_pattern = {96{1'b0}};correction_pattern[51]=1'b1;
			end
			8'b01001100: begin
				correction_pattern = {96{1'b0}};correction_pattern[52]=1'b1;
			end
			8'b00001110: begin
				correction_pattern = {96{1'b0}};correction_pattern[53]=1'b1;
			end
			8'b00010011: begin
				correction_pattern = {96{1'b0}};correction_pattern[54]=1'b1;
			end
			8'b11100000: begin
				correction_pattern = {96{1'b0}};correction_pattern[55]=1'b1;
			end
			8'b11100011: begin
				correction_pattern = {96{1'b0}};correction_pattern[56]=1'b1;
			end
			8'b01111100: begin
				correction_pattern = {96{1'b0}};correction_pattern[57]=1'b1;
			end
			8'b10011110: begin
				correction_pattern = {96{1'b0}};correction_pattern[58]=1'b1;
			end
			8'b10011101: begin
				correction_pattern = {96{1'b0}};correction_pattern[59]=1'b1;
			end
			8'b01110011: begin
				correction_pattern = {96{1'b0}};correction_pattern[60]=1'b1;
			end
			8'b01100111: begin
				correction_pattern = {96{1'b0}};correction_pattern[61]=1'b1;
			end
			8'b11001011: begin
				correction_pattern = {96{1'b0}};correction_pattern[62]=1'b1;
			end
			8'b10111100: begin
				correction_pattern = {96{1'b0}};correction_pattern[63]=1'b1;
			end
			8'b10101101: begin
				correction_pattern = {96{1'b0}};correction_pattern[64]=1'b1;
			end
			8'b11011010: begin
				correction_pattern = {96{1'b0}};correction_pattern[65]=1'b1;
			end
			8'b01110110: begin
				correction_pattern = {96{1'b0}};correction_pattern[66]=1'b1;
			end
			8'b01010111: begin
				correction_pattern = {96{1'b0}};correction_pattern[67]=1'b1;
			end
			8'b10111001: begin
				correction_pattern = {96{1'b0}};correction_pattern[68]=1'b1;
			end
			8'b10101011: begin
				correction_pattern = {96{1'b0}};correction_pattern[69]=1'b1;
			end
			8'b01101101: begin
				correction_pattern = {96{1'b0}};correction_pattern[70]=1'b1;
			end
			8'b11010110: begin
				correction_pattern = {96{1'b0}};correction_pattern[71]=1'b1;
			end
			8'b11000111: begin
				correction_pattern = {96{1'b0}};correction_pattern[72]=1'b1;
			end
			8'b11111000: begin
				correction_pattern = {96{1'b0}};correction_pattern[73]=1'b1;
			end
			8'b00111110: begin
				correction_pattern = {96{1'b0}};correction_pattern[74]=1'b1;
			end
			8'b00111101: begin
				correction_pattern = {96{1'b0}};correction_pattern[75]=1'b1;
			end
			8'b11010011: begin
				correction_pattern = {96{1'b0}};correction_pattern[76]=1'b1;
			end
			8'b01101011: begin
				correction_pattern = {96{1'b0}};correction_pattern[77]=1'b1;
			end
			8'b10100111: begin
				correction_pattern = {96{1'b0}};correction_pattern[78]=1'b1;
			end
			8'b11011100: begin
				correction_pattern = {96{1'b0}};correction_pattern[79]=1'b1;
			end
			8'b11001101: begin
				correction_pattern = {96{1'b0}};correction_pattern[80]=1'b1;
			end
			8'b10110110: begin
				correction_pattern = {96{1'b0}};correction_pattern[81]=1'b1;
			end
			8'b01111010: begin
				correction_pattern = {96{1'b0}};correction_pattern[82]=1'b1;
			end
			8'b00111011: begin
				correction_pattern = {96{1'b0}};correction_pattern[83]=1'b1;
			end
			8'b11010101: begin
				correction_pattern = {96{1'b0}};correction_pattern[84]=1'b1;
			end
			8'b11100101: begin
				correction_pattern = {96{1'b0}};correction_pattern[85]=1'b1;
			end
			8'b01001111: begin
				correction_pattern = {96{1'b0}};correction_pattern[86]=1'b1;
			end
			8'b10111010: begin
				correction_pattern = {96{1'b0}};correction_pattern[87]=1'b1;
			end
			8'b11101010: begin
				correction_pattern = {96{1'b0}};correction_pattern[88]=1'b1;
			end
			8'b00011111: begin
				correction_pattern = {96{1'b0}};correction_pattern[89]=1'b1;
			end
			8'b10110101: begin
				correction_pattern = {96{1'b0}};correction_pattern[90]=1'b1;
			end
			8'b01110101: begin
				correction_pattern = {96{1'b0}};correction_pattern[91]=1'b1;
			end
			8'b11001110: begin
				correction_pattern = {96{1'b0}};correction_pattern[92]=1'b1;
			end
			8'b11110010: begin
				correction_pattern = {96{1'b0}};correction_pattern[93]=1'b1;
			end
			8'b11011001: begin
				correction_pattern = {96{1'b0}};correction_pattern[94]=1'b1;
			end
			8'b00101111: begin
				correction_pattern = {96{1'b0}};correction_pattern[95]=1'b1;
			end
			8'b00000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b01000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b10000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_104_96_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [8-1:0] stored_data_edc = extended_hamming_code_104_96_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [96-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_104_96_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_128_min_width (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_136_128_f
//Compute 8 bits Error Detection Code from a 128 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used 2 times (syndrom bits 0 1)
//  input bit   1 used 2 times (syndrom bits 2 3)
//  input bit   2 used 2 times (syndrom bits 4 5)
//  input bit   3 used 2 times (syndrom bits 6 7)
//  input bit   4 used 2 times (syndrom bits 4 6)
//  input bit   5 used 2 times (syndrom bits 5 7)
//  input bit   6 used 2 times (syndrom bits 0 2)
//  input bit   7 used 2 times (syndrom bits 1 3)
//  input bit   8 used 2 times (syndrom bits 0 3)
//  input bit   9 used 2 times (syndrom bits 1 2)
//  input bit  10 used 2 times (syndrom bits 4 7)
//  input bit  11 used 2 times (syndrom bits 5 6)
//  input bit  12 used 2 times (syndrom bits 1 5)
//  input bit  13 used 2 times (syndrom bits 2 6)
//  input bit  14 used 2 times (syndrom bits 3 7)
//  input bit  15 used 2 times (syndrom bits 0 4)
//  input bit  16 used 2 times (syndrom bits 3 4)
//  input bit  17 used 2 times (syndrom bits 0 7)
//  input bit  18 used 2 times (syndrom bits 1 6)
//  input bit  19 used 2 times (syndrom bits 2 5)
//  input bit  20 used 2 times (syndrom bits 2 7)
//  input bit  21 used 2 times (syndrom bits 0 5)
//  input bit  22 used 2 times (syndrom bits 3 6)
//  input bit  23 used 2 times (syndrom bits 1 4)
//  input bit  24 used 2 times (syndrom bits 1 7)
//  input bit  25 used 2 times (syndrom bits 2 4)
//  input bit  26 used 2 times (syndrom bits 0 6)
//  input bit  27 used 2 times (syndrom bits 3 5)
//  input bit  28 used 3 times (syndrom bits 3 5 6)
//  input bit  29 used 3 times (syndrom bits 0 2 4)
//  input bit  30 used 3 times (syndrom bits 0 1 7)
//  input bit  31 used 3 times (syndrom bits 1 4 7)
//  input bit  32 used 3 times (syndrom bits 2 3 5)
//  input bit  33 used 3 times (syndrom bits 2 3 6)
//  input bit  34 used 3 times (syndrom bits 1 5 6)
//  input bit  35 used 3 times (syndrom bits 0 4 7)
//  input bit  36 used 3 times (syndrom bits 4 6 7)
//  input bit  37 used 3 times (syndrom bits 0 1 5)
//  input bit  38 used 3 times (syndrom bits 0 2 3)
//  input bit  39 used 3 times (syndrom bits 1 2 3)
//  input bit  40 used 3 times (syndrom bits 4 5 7)
//  input bit  41 used 3 times (syndrom bits 5 6 7)
//  input bit  42 used 3 times (syndrom bits 2 4 6)
//  input bit  43 used 3 times (syndrom bits 0 1 3)
//  input bit  44 used 3 times (syndrom bits 1 3 6)
//  input bit  45 used 3 times (syndrom bits 0 4 5)
//  input bit  46 used 3 times (syndrom bits 0 2 7)
//  input bit  47 used 3 times (syndrom bits 2 4 7)
//  input bit  48 used 3 times (syndrom bits 1 3 5)
//  input bit  49 used 3 times (syndrom bits 2 5 6)
//  input bit  50 used 3 times (syndrom bits 3 6 7)
//  input bit  51 used 3 times (syndrom bits 0 1 4)
//  input bit  52 used 3 times (syndrom bits 1 4 6)
//  input bit  53 used 3 times (syndrom bits 0 3 7)
//  input bit  54 used 3 times (syndrom bits 0 2 5)
//  input bit  55 used 3 times (syndrom bits 2 5 7)
//  input bit  56 used 3 times (syndrom bits 1 3 4)
//  input bit  57 used 3 times (syndrom bits 3 4 6)
//  input bit  58 used 3 times (syndrom bits 1 2 6)
//  input bit  59 used 3 times (syndrom bits 0 5 7)
//  input bit  60 used 3 times (syndrom bits 1 5 7)
//  input bit  61 used 3 times (syndrom bits 0 2 6)
//  input bit  62 used 3 times (syndrom bits 0 3 4)
//  input bit  63 used 3 times (syndrom bits 2 3 4)
//  input bit  64 used 3 times (syndrom bits 4 5 6)
//  input bit  65 used 3 times (syndrom bits 1 6 7)
//  input bit  66 used 3 times (syndrom bits 1 3 7)
//  input bit  67 used 3 times (syndrom bits 1 2 5)
//  input bit  68 used 3 times (syndrom bits 0 3 5)
//  input bit  69 used 3 times (syndrom bits 0 1 2)
//  input bit  70 used 3 times (syndrom bits 0 6 7)
//  input bit  71 used 3 times (syndrom bits 3 4 7)
//  input bit  72 used 3 times (syndrom bits 0 4 6)
//  input bit  73 used 3 times (syndrom bits 2 4 5)
//  input bit  74 used 3 times (syndrom bits 2 6 7)
//  input bit  75 used 3 times (syndrom bits 3 5 7)
//  input bit  76 used 3 times (syndrom bits 1 4 5)
//  input bit  77 used 3 times (syndrom bits 1 2 4)
//  input bit  78 used 3 times (syndrom bits 0 3 6)
//  input bit  79 used 3 times (syndrom bits 2 3 7)
//  input bit  80 used 3 times (syndrom bits 0 1 6)
//  input bit  81 used 3 times (syndrom bits 0 5 6)
//  input bit  82 used 3 times (syndrom bits 3 4 5)
//  input bit  83 used 3 times (syndrom bits 1 2 7)
//  input bit  84 used 4 times (syndrom bits 1 2 5 7)
//  input bit  85 used 4 times (syndrom bits 0 3 4 6)
//  input bit  86 used 4 times (syndrom bits 1 3 4 6)
//  input bit  87 used 4 times (syndrom bits 0 2 5 7)
//  input bit  88 used 4 times (syndrom bits 0 2 3 7)
//  input bit  89 used 4 times (syndrom bits 1 4 5 6)
//  input bit  90 used 4 times (syndrom bits 0 4 5 6)
//  input bit  91 used 4 times (syndrom bits 1 2 3 7)
//  input bit  92 used 4 times (syndrom bits 1 2 4 7)
//  input bit  93 used 4 times (syndrom bits 0 3 5 6)
//  input bit  94 used 4 times (syndrom bits 1 3 5 6)
//  input bit  95 used 4 times (syndrom bits 0 2 4 7)
//  input bit  96 used 4 times (syndrom bits 0 2 6 7)
//  input bit  97 used 4 times (syndrom bits 1 3 4 5)
//  input bit  98 used 4 times (syndrom bits 0 3 4 5)
//  input bit  99 used 4 times (syndrom bits 1 2 6 7)
//  input bit 100 used 4 times (syndrom bits 0 1 2 7)
//  input bit 101 used 4 times (syndrom bits 3 4 5 6)
//  input bit 102 used 4 times (syndrom bits 2 3 4 6)
//  input bit 103 used 4 times (syndrom bits 0 1 5 7)
//  input bit 104 used 4 times (syndrom bits 1 5 6 7)
//  input bit 105 used 4 times (syndrom bits 0 2 3 4)
//  input bit 106 used 4 times (syndrom bits 0 1 3 4)
//  input bit 107 used 4 times (syndrom bits 2 5 6 7)
//  input bit 108 used 4 times (syndrom bits 2 4 5 7)
//  input bit 109 used 4 times (syndrom bits 0 1 3 6)
//  input bit 110 used 4 times (syndrom bits 0 2 3 6)
//  input bit 111 used 4 times (syndrom bits 1 4 5 7)
//  input bit 112 used 4 times (syndrom bits 1 3 5 7)
//  input bit 113 used 4 times (syndrom bits 0 2 4 6)
//  input bit 114 used 4 times (syndrom bits 0 1 4 6)
//  input bit 115 used 4 times (syndrom bits 2 3 5 7)
//  input bit 116 used 4 times (syndrom bits 2 3 4 5)
//  input bit 117 used 4 times (syndrom bits 0 1 6 7)
//  input bit 118 used 4 times (syndrom bits 0 5 6 7)
//  input bit 119 used 4 times (syndrom bits 1 2 3 4)
//  input bit 120 used 4 times (syndrom bits 1 2 3 6)
//  input bit 121 used 4 times (syndrom bits 0 4 5 7)
//  input bit 122 used 4 times (syndrom bits 0 1 4 7)
//  input bit 123 used 4 times (syndrom bits 2 3 5 6)
//  input bit 124 used 4 times (syndrom bits 0 2 3 5)
//  input bit 125 used 4 times (syndrom bits 1 4 6 7)
//  input bit 126 used 4 times (syndrom bits 4 5 6 7)
//  input bit 127 used 4 times (syndrom bits 0 1 2 3)
function [8-1:0] hamming_code_136_128_f;
    input [128-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[  0]^in[  6]^in[  8]^in[ 15]^in[ 17]^in[ 21]^in[ 26]^in[ 29]^in[ 30]^in[ 35]^in[ 37]^in[ 38]^in[ 43]^in[ 45]^in[ 46]^in[ 51]^in[ 53]^in[ 54]^in[ 59]^in[ 61]^in[ 62]^in[ 68]^in[ 69]^in[ 70]^in[ 72]^in[ 78]^in[ 80]^in[ 81]^in[ 85]^in[ 87]^in[ 88]^in[ 90]^in[ 93]^in[ 95]^in[ 96]^in[ 98]^in[100]^in[103]^in[105]^in[106]^in[109]^in[110]^in[113]^in[114]^in[117]^in[118]^in[121]^in[122]^in[124]^in[127];//50 inputs
        syndrom[1] = in[  0]^in[  7]^in[  9]^in[ 12]^in[ 18]^in[ 23]^in[ 24]^in[ 30]^in[ 31]^in[ 34]^in[ 37]^in[ 39]^in[ 43]^in[ 44]^in[ 48]^in[ 51]^in[ 52]^in[ 56]^in[ 58]^in[ 60]^in[ 65]^in[ 66]^in[ 67]^in[ 69]^in[ 76]^in[ 77]^in[ 80]^in[ 83]^in[ 84]^in[ 86]^in[ 89]^in[ 91]^in[ 92]^in[ 94]^in[ 97]^in[ 99]^in[100]^in[103]^in[104]^in[106]^in[109]^in[111]^in[112]^in[114]^in[117]^in[119]^in[120]^in[122]^in[125]^in[127];//50 inputs
        syndrom[2] = in[  1]^in[  6]^in[  9]^in[ 13]^in[ 19]^in[ 20]^in[ 25]^in[ 29]^in[ 32]^in[ 33]^in[ 38]^in[ 39]^in[ 42]^in[ 46]^in[ 47]^in[ 49]^in[ 54]^in[ 55]^in[ 58]^in[ 61]^in[ 63]^in[ 67]^in[ 69]^in[ 73]^in[ 74]^in[ 77]^in[ 79]^in[ 83]^in[ 84]^in[ 87]^in[ 88]^in[ 91]^in[ 92]^in[ 95]^in[ 96]^in[ 99]^in[100]^in[102]^in[105]^in[107]^in[108]^in[110]^in[113]^in[115]^in[116]^in[119]^in[120]^in[123]^in[124]^in[127];//50 inputs
        syndrom[3] = in[  1]^in[  7]^in[  8]^in[ 14]^in[ 16]^in[ 22]^in[ 27]^in[ 28]^in[ 32]^in[ 33]^in[ 38]^in[ 39]^in[ 43]^in[ 44]^in[ 48]^in[ 50]^in[ 53]^in[ 56]^in[ 57]^in[ 62]^in[ 63]^in[ 66]^in[ 68]^in[ 71]^in[ 75]^in[ 78]^in[ 79]^in[ 82]^in[ 85]^in[ 86]^in[ 88]^in[ 91]^in[ 93]^in[ 94]^in[ 97]^in[ 98]^in[101]^in[102]^in[105]^in[106]^in[109]^in[110]^in[112]^in[115]^in[116]^in[119]^in[120]^in[123]^in[124]^in[127];//50 inputs
        syndrom[4] = in[  2]^in[  4]^in[ 10]^in[ 15]^in[ 16]^in[ 23]^in[ 25]^in[ 29]^in[ 31]^in[ 35]^in[ 36]^in[ 40]^in[ 42]^in[ 45]^in[ 47]^in[ 51]^in[ 52]^in[ 56]^in[ 57]^in[ 62]^in[ 63]^in[ 64]^in[ 71]^in[ 72]^in[ 73]^in[ 76]^in[ 77]^in[ 82]^in[ 85]^in[ 86]^in[ 89]^in[ 90]^in[ 92]^in[ 95]^in[ 97]^in[ 98]^in[101]^in[102]^in[105]^in[106]^in[108]^in[111]^in[113]^in[114]^in[116]^in[119]^in[121]^in[122]^in[125]^in[126];//50 inputs
        syndrom[5] = in[  2]^in[  5]^in[ 11]^in[ 12]^in[ 19]^in[ 21]^in[ 27]^in[ 28]^in[ 32]^in[ 34]^in[ 37]^in[ 40]^in[ 41]^in[ 45]^in[ 48]^in[ 49]^in[ 54]^in[ 55]^in[ 59]^in[ 60]^in[ 64]^in[ 67]^in[ 68]^in[ 73]^in[ 75]^in[ 76]^in[ 81]^in[ 82]^in[ 84]^in[ 87]^in[ 89]^in[ 90]^in[ 93]^in[ 94]^in[ 97]^in[ 98]^in[101]^in[103]^in[104]^in[107]^in[108]^in[111]^in[112]^in[115]^in[116]^in[118]^in[121]^in[123]^in[124]^in[126];//50 inputs
        syndrom[6] = in[  3]^in[  4]^in[ 11]^in[ 13]^in[ 18]^in[ 22]^in[ 26]^in[ 28]^in[ 33]^in[ 34]^in[ 36]^in[ 41]^in[ 42]^in[ 44]^in[ 49]^in[ 50]^in[ 52]^in[ 57]^in[ 58]^in[ 61]^in[ 64]^in[ 65]^in[ 70]^in[ 72]^in[ 74]^in[ 78]^in[ 80]^in[ 81]^in[ 85]^in[ 86]^in[ 89]^in[ 90]^in[ 93]^in[ 94]^in[ 96]^in[ 99]^in[101]^in[102]^in[104]^in[107]^in[109]^in[110]^in[113]^in[114]^in[117]^in[118]^in[120]^in[123]^in[125]^in[126];//50 inputs
        syndrom[7] = in[  3]^in[  5]^in[ 10]^in[ 14]^in[ 17]^in[ 20]^in[ 24]^in[ 30]^in[ 31]^in[ 35]^in[ 36]^in[ 40]^in[ 41]^in[ 46]^in[ 47]^in[ 50]^in[ 53]^in[ 55]^in[ 59]^in[ 60]^in[ 65]^in[ 66]^in[ 70]^in[ 71]^in[ 74]^in[ 75]^in[ 79]^in[ 83]^in[ 84]^in[ 87]^in[ 88]^in[ 91]^in[ 92]^in[ 95]^in[ 96]^in[ 99]^in[100]^in[103]^in[104]^in[107]^in[108]^in[111]^in[112]^in[115]^in[117]^in[118]^in[121]^in[122]^in[125]^in[126];//50 inputs
        hamming_code_136_128_f = syndrom;
    end
endfunction
wire [8-1:0] stored_data_edc = hamming_code_136_128_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_128_min_width (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [9-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [9-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_137_128_f
//Compute 9 bits Error Detection Code from a 128 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used 3 times (syndrom bits 0 1 2)
//  input bit   1 used 3 times (syndrom bits 3 4 5)
//  input bit   2 used 3 times (syndrom bits 6 7 8)
//  input bit   3 used 3 times (syndrom bits 3 6 7)
//  input bit   4 used 3 times (syndrom bits 4 5 8)
//  input bit   5 used 3 times (syndrom bits 0 1 8)
//  input bit   6 used 3 times (syndrom bits 0 2 4)
//  input bit   7 used 3 times (syndrom bits 1 2 5)
//  input bit   8 used 3 times (syndrom bits 2 6 7)
//  input bit   9 used 3 times (syndrom bits 1 3 6)
//  input bit  10 used 3 times (syndrom bits 3 5 7)
//  input bit  11 used 3 times (syndrom bits 0 4 8)
//  input bit  12 used 3 times (syndrom bits 0 3 4)
//  input bit  13 used 3 times (syndrom bits 5 7 8)
//  input bit  14 used 3 times (syndrom bits 1 2 6)
//  input bit  15 used 3 times (syndrom bits 1 6 8)
//  input bit  16 used 3 times (syndrom bits 2 5 7)
//  input bit  17 used 3 times (syndrom bits 0 4 7)
//  input bit  18 used 3 times (syndrom bits 0 2 3)
//  input bit  19 used 3 times (syndrom bits 3 4 6)
//  input bit  20 used 3 times (syndrom bits 1 5 8)
//  input bit  21 used 3 times (syndrom bits 1 3 5)
//  input bit  22 used 3 times (syndrom bits 4 6 8)
//  input bit  23 used 3 times (syndrom bits 0 2 7)
//  input bit  24 used 3 times (syndrom bits 0 2 8)
//  input bit  25 used 3 times (syndrom bits 4 6 7)
//  input bit  26 used 3 times (syndrom bits 1 5 7)
//  input bit  27 used 3 times (syndrom bits 3 5 6)
//  input bit  28 used 3 times (syndrom bits 1 3 4)
//  input bit  29 used 3 times (syndrom bits 0 2 5)
//  input bit  30 used 3 times (syndrom bits 0 3 8)
//  input bit  31 used 3 times (syndrom bits 1 2 8)
//  input bit  32 used 3 times (syndrom bits 2 4 6)
//  input bit  33 used 3 times (syndrom bits 4 7 8)
//  input bit  34 used 3 times (syndrom bits 1 6 7)
//  input bit  35 used 3 times (syndrom bits 0 3 5)
//  input bit  36 used 3 times (syndrom bits 0 3 7)
//  input bit  37 used 3 times (syndrom bits 1 5 6)
//  input bit  38 used 3 times (syndrom bits 2 4 8)
//  input bit  39 used 3 times (syndrom bits 1 4 8)
//  input bit  40 used 3 times (syndrom bits 2 5 6)
//  input bit  41 used 3 times (syndrom bits 0 3 6)
//  input bit  42 used 3 times (syndrom bits 0 5 7)
//  input bit  43 used 3 times (syndrom bits 2 3 7)
//  input bit  44 used 3 times (syndrom bits 3 4 8)
//  input bit  45 used 3 times (syndrom bits 1 4 7)
//  input bit  46 used 3 times (syndrom bits 1 7 8)
//  input bit  47 used 3 times (syndrom bits 0 2 6)
//  input bit  48 used 3 times (syndrom bits 2 5 8)
//  input bit  49 used 3 times (syndrom bits 0 5 6)
//  input bit  50 used 3 times (syndrom bits 1 4 5)
//  input bit  51 used 3 times (syndrom bits 0 1 3)
//  input bit  52 used 3 times (syndrom bits 2 3 4)
//  input bit  53 used 3 times (syndrom bits 3 6 8)
//  input bit  54 used 3 times (syndrom bits 0 6 7)
//  input bit  55 used 3 times (syndrom bits 2 7 8)
//  input bit  56 used 3 times (syndrom bits 1 2 4)
//  input bit  57 used 3 times (syndrom bits 4 5 7)
//  input bit  58 used 3 times (syndrom bits 0 1 5)
//  input bit  59 used 3 times (syndrom bits 5 6 8)
//  input bit  60 used 3 times (syndrom bits 1 3 8)
//  input bit  61 used 3 times (syndrom bits 2 3 6)
//  input bit  62 used 3 times (syndrom bits 0 4 6)
//  input bit  63 used 3 times (syndrom bits 0 7 8)
//  input bit  64 used 3 times (syndrom bits 3 4 7)
//  input bit  65 used 3 times (syndrom bits 1 2 7)
//  input bit  66 used 3 times (syndrom bits 2 4 5)
//  input bit  67 used 3 times (syndrom bits 3 5 8)
//  input bit  68 used 3 times (syndrom bits 0 1 6)
//  input bit  69 used 3 times (syndrom bits 0 1 4)
//  input bit  70 used 3 times (syndrom bits 5 6 7)
//  input bit  71 used 3 times (syndrom bits 2 3 8)
//  input bit  72 used 3 times (syndrom bits 3 7 8)
//  input bit  73 used 3 times (syndrom bits 2 6 8)
//  input bit  74 used 3 times (syndrom bits 0 4 5)
//  input bit  75 used 3 times (syndrom bits 0 1 7)
//  input bit  76 used 3 times (syndrom bits 1 4 6)
//  input bit  77 used 3 times (syndrom bits 2 3 5)
//  input bit  78 used 3 times (syndrom bits 4 5 6)
//  input bit  79 used 3 times (syndrom bits 1 2 3)
//  input bit  80 used 3 times (syndrom bits 0 5 8)
//  input bit  81 used 3 times (syndrom bits 2 4 7)
//  input bit  82 used 3 times (syndrom bits 1 3 7)
//  input bit  83 used 3 times (syndrom bits 0 6 8)
//  input bit  84 used 5 times (syndrom bits 0 3 6 7 8)
//  input bit  85 used 5 times (syndrom bits 0 1 2 4 5)
//  input bit  86 used 5 times (syndrom bits 1 2 4 5 8)
//  input bit  87 used 5 times (syndrom bits 1 2 3 6 7)
//  input bit  88 used 5 times (syndrom bits 3 4 5 6 7)
//  input bit  89 used 5 times (syndrom bits 0 4 6 7 8)
//  input bit  90 used 5 times (syndrom bits 0 1 3 5 8)
//  input bit  91 used 5 times (syndrom bits 0 2 3 5 8)
//  input bit  92 used 5 times (syndrom bits 1 2 4 6 7)
//  input bit  93 used 5 times (syndrom bits 1 2 6 7 8)
//  input bit  94 used 5 times (syndrom bits 0 2 3 4 5)
//  input bit  95 used 5 times (syndrom bits 0 1 3 4 5)
//  input bit  96 used 5 times (syndrom bits 3 4 6 7 8)
//  input bit  97 used 5 times (syndrom bits 0 5 6 7 8)
//  input bit  98 used 5 times (syndrom bits 0 1 2 6 7)
//  input bit  99 used 5 times (syndrom bits 1 2 3 5 8)
//  input bit 100 used 5 times (syndrom bits 1 2 3 4 8)
//  input bit 101 used 5 times (syndrom bits 0 4 5 6 7)
//  input bit 102 used 5 times (syndrom bits 1 4 5 6 7)
//  input bit 103 used 5 times (syndrom bits 0 2 3 4 8)
//  input bit 104 used 5 times (syndrom bits 0 2 3 6 8)
//  input bit 105 used 5 times (syndrom bits 0 1 2 5 7)
//  input bit 106 used 5 times (syndrom bits 1 3 5 7 8)
//  input bit 107 used 5 times (syndrom bits 4 5 6 7 8)
//  input bit 108 used 5 times (syndrom bits 0 1 3 4 6)
//  input bit 109 used 5 times (syndrom bits 1 2 3 4 6)
//  input bit 110 used 5 times (syndrom bits 0 2 5 7 8)
//  input bit 111 used 5 times (syndrom bits 0 2 5 6 7)
//  input bit 112 used 5 times (syndrom bits 0 1 3 4 8)
//  input bit 113 used 5 times (syndrom bits 1 3 4 5 8)
//  input bit 114 used 5 times (syndrom bits 2 4 6 7 8)
//  input bit 115 used 5 times (syndrom bits 1 2 5 6 7)
//  input bit 116 used 5 times (syndrom bits 0 2 3 6 7)
//  input bit 117 used 5 times (syndrom bits 0 1 2 3 5)
//  input bit 118 used 5 times (syndrom bits 0 3 4 5 8)
//  input bit 119 used 5 times (syndrom bits 1 4 6 7 8)
//  input bit 120 used 5 times (syndrom bits 1 3 4 7 8)
//  input bit 121 used 5 times (syndrom bits 0 2 5 6 8)
//  input bit 122 used 5 times (syndrom bits 0 2 4 5 6)
//  input bit 123 used 5 times (syndrom bits 0 1 3 6 7)
//  input bit 124 used 5 times (syndrom bits 1 2 3 5 7)
//  input bit 125 used 5 times (syndrom bits 1 4 5 7 8)
//  input bit 126 used 5 times (syndrom bits 2 3 4 6 8)
//  input bit 127 used 5 times (syndrom bits 0 3 4 6 8)
function [9-1:0] extended_hamming_code_137_128_f;
    input [128-1:0] in;
    reg [9-1:0] syndrom;
    begin
        syndrom[0] = in[  0]^in[  5]^in[  6]^in[ 11]^in[ 12]^in[ 17]^in[ 18]^in[ 23]^in[ 24]^in[ 29]^in[ 30]^in[ 35]^in[ 36]^in[ 41]^in[ 42]^in[ 47]^in[ 49]^in[ 51]^in[ 54]^in[ 58]^in[ 62]^in[ 63]^in[ 68]^in[ 69]^in[ 74]^in[ 75]^in[ 80]^in[ 83]^in[ 84]^in[ 85]^in[ 89]^in[ 90]^in[ 91]^in[ 94]^in[ 95]^in[ 97]^in[ 98]^in[101]^in[103]^in[104]^in[105]^in[108]^in[110]^in[111]^in[112]^in[116]^in[117]^in[118]^in[121]^in[122]^in[123]^in[127];//52 inputs
        syndrom[1] = in[  0]^in[  5]^in[  7]^in[  9]^in[ 14]^in[ 15]^in[ 20]^in[ 21]^in[ 26]^in[ 28]^in[ 31]^in[ 34]^in[ 37]^in[ 39]^in[ 45]^in[ 46]^in[ 50]^in[ 51]^in[ 56]^in[ 58]^in[ 60]^in[ 65]^in[ 68]^in[ 69]^in[ 75]^in[ 76]^in[ 79]^in[ 82]^in[ 85]^in[ 86]^in[ 87]^in[ 90]^in[ 92]^in[ 93]^in[ 95]^in[ 98]^in[ 99]^in[100]^in[102]^in[105]^in[106]^in[108]^in[109]^in[112]^in[113]^in[115]^in[117]^in[119]^in[120]^in[123]^in[124]^in[125];//52 inputs
        syndrom[2] = in[  0]^in[  6]^in[  7]^in[  8]^in[ 14]^in[ 16]^in[ 18]^in[ 23]^in[ 24]^in[ 29]^in[ 31]^in[ 32]^in[ 38]^in[ 40]^in[ 43]^in[ 47]^in[ 48]^in[ 52]^in[ 55]^in[ 56]^in[ 61]^in[ 65]^in[ 66]^in[ 71]^in[ 73]^in[ 77]^in[ 79]^in[ 81]^in[ 85]^in[ 86]^in[ 87]^in[ 91]^in[ 92]^in[ 93]^in[ 94]^in[ 98]^in[ 99]^in[100]^in[103]^in[104]^in[105]^in[109]^in[110]^in[111]^in[114]^in[115]^in[116]^in[117]^in[121]^in[122]^in[124]^in[126];//52 inputs
        syndrom[3] = in[  1]^in[  3]^in[  9]^in[ 10]^in[ 12]^in[ 18]^in[ 19]^in[ 21]^in[ 27]^in[ 28]^in[ 30]^in[ 35]^in[ 36]^in[ 41]^in[ 43]^in[ 44]^in[ 51]^in[ 52]^in[ 53]^in[ 60]^in[ 61]^in[ 64]^in[ 67]^in[ 71]^in[ 72]^in[ 77]^in[ 79]^in[ 82]^in[ 84]^in[ 87]^in[ 88]^in[ 90]^in[ 91]^in[ 94]^in[ 95]^in[ 96]^in[ 99]^in[100]^in[103]^in[104]^in[106]^in[108]^in[109]^in[112]^in[113]^in[116]^in[117]^in[118]^in[120]^in[123]^in[124]^in[126]^in[127];//53 inputs
        syndrom[4] = in[  1]^in[  4]^in[  6]^in[ 11]^in[ 12]^in[ 17]^in[ 19]^in[ 22]^in[ 25]^in[ 28]^in[ 32]^in[ 33]^in[ 38]^in[ 39]^in[ 44]^in[ 45]^in[ 50]^in[ 52]^in[ 56]^in[ 57]^in[ 62]^in[ 64]^in[ 66]^in[ 69]^in[ 74]^in[ 76]^in[ 78]^in[ 81]^in[ 85]^in[ 86]^in[ 88]^in[ 89]^in[ 92]^in[ 94]^in[ 95]^in[ 96]^in[100]^in[101]^in[102]^in[103]^in[107]^in[108]^in[109]^in[112]^in[113]^in[114]^in[118]^in[119]^in[120]^in[122]^in[125]^in[126]^in[127];//53 inputs
        syndrom[5] = in[  1]^in[  4]^in[  7]^in[ 10]^in[ 13]^in[ 16]^in[ 20]^in[ 21]^in[ 26]^in[ 27]^in[ 29]^in[ 35]^in[ 37]^in[ 40]^in[ 42]^in[ 48]^in[ 49]^in[ 50]^in[ 57]^in[ 58]^in[ 59]^in[ 66]^in[ 67]^in[ 70]^in[ 74]^in[ 77]^in[ 78]^in[ 80]^in[ 85]^in[ 86]^in[ 88]^in[ 90]^in[ 91]^in[ 94]^in[ 95]^in[ 97]^in[ 99]^in[101]^in[102]^in[105]^in[106]^in[107]^in[110]^in[111]^in[113]^in[115]^in[117]^in[118]^in[121]^in[122]^in[124]^in[125];//52 inputs
        syndrom[6] = in[  2]^in[  3]^in[  8]^in[  9]^in[ 14]^in[ 15]^in[ 19]^in[ 22]^in[ 25]^in[ 27]^in[ 32]^in[ 34]^in[ 37]^in[ 40]^in[ 41]^in[ 47]^in[ 49]^in[ 53]^in[ 54]^in[ 59]^in[ 61]^in[ 62]^in[ 68]^in[ 70]^in[ 73]^in[ 76]^in[ 78]^in[ 83]^in[ 84]^in[ 87]^in[ 88]^in[ 89]^in[ 92]^in[ 93]^in[ 96]^in[ 97]^in[ 98]^in[101]^in[102]^in[104]^in[107]^in[108]^in[109]^in[111]^in[114]^in[115]^in[116]^in[119]^in[121]^in[122]^in[123]^in[126]^in[127];//53 inputs
        syndrom[7] = in[  2]^in[  3]^in[  8]^in[ 10]^in[ 13]^in[ 16]^in[ 17]^in[ 23]^in[ 25]^in[ 26]^in[ 33]^in[ 34]^in[ 36]^in[ 42]^in[ 43]^in[ 45]^in[ 46]^in[ 54]^in[ 55]^in[ 57]^in[ 63]^in[ 64]^in[ 65]^in[ 70]^in[ 72]^in[ 75]^in[ 81]^in[ 82]^in[ 84]^in[ 87]^in[ 88]^in[ 89]^in[ 92]^in[ 93]^in[ 96]^in[ 97]^in[ 98]^in[101]^in[102]^in[105]^in[106]^in[107]^in[110]^in[111]^in[114]^in[115]^in[116]^in[119]^in[120]^in[123]^in[124]^in[125];//52 inputs
        syndrom[8] = in[  2]^in[  4]^in[  5]^in[ 11]^in[ 13]^in[ 15]^in[ 20]^in[ 22]^in[ 24]^in[ 30]^in[ 31]^in[ 33]^in[ 38]^in[ 39]^in[ 44]^in[ 46]^in[ 48]^in[ 53]^in[ 55]^in[ 59]^in[ 60]^in[ 63]^in[ 67]^in[ 71]^in[ 72]^in[ 73]^in[ 80]^in[ 83]^in[ 84]^in[ 86]^in[ 89]^in[ 90]^in[ 91]^in[ 93]^in[ 96]^in[ 97]^in[ 99]^in[100]^in[103]^in[104]^in[106]^in[107]^in[110]^in[112]^in[113]^in[114]^in[118]^in[119]^in[120]^in[121]^in[125]^in[126]^in[127];//53 inputs
        extended_hamming_code_137_128_f = syndrom;
    end
endfunction
wire [9-1:0] stored_data_edc = extended_hamming_code_137_128_f(i_stored_data);
wire [9-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_128_min_width (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [9-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [9-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [128-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_137_128_f
//Compute 9 bits Error Detection Code from a 128 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used 3 times (syndrom bits 0 1 2)
//  input bit   1 used 3 times (syndrom bits 3 4 5)
//  input bit   2 used 3 times (syndrom bits 6 7 8)
//  input bit   3 used 3 times (syndrom bits 3 6 7)
//  input bit   4 used 3 times (syndrom bits 4 5 8)
//  input bit   5 used 3 times (syndrom bits 0 1 8)
//  input bit   6 used 3 times (syndrom bits 0 2 4)
//  input bit   7 used 3 times (syndrom bits 1 2 5)
//  input bit   8 used 3 times (syndrom bits 2 6 7)
//  input bit   9 used 3 times (syndrom bits 1 3 6)
//  input bit  10 used 3 times (syndrom bits 3 5 7)
//  input bit  11 used 3 times (syndrom bits 0 4 8)
//  input bit  12 used 3 times (syndrom bits 0 3 4)
//  input bit  13 used 3 times (syndrom bits 5 7 8)
//  input bit  14 used 3 times (syndrom bits 1 2 6)
//  input bit  15 used 3 times (syndrom bits 1 6 8)
//  input bit  16 used 3 times (syndrom bits 2 5 7)
//  input bit  17 used 3 times (syndrom bits 0 4 7)
//  input bit  18 used 3 times (syndrom bits 0 2 3)
//  input bit  19 used 3 times (syndrom bits 3 4 6)
//  input bit  20 used 3 times (syndrom bits 1 5 8)
//  input bit  21 used 3 times (syndrom bits 1 3 5)
//  input bit  22 used 3 times (syndrom bits 4 6 8)
//  input bit  23 used 3 times (syndrom bits 0 2 7)
//  input bit  24 used 3 times (syndrom bits 0 2 8)
//  input bit  25 used 3 times (syndrom bits 4 6 7)
//  input bit  26 used 3 times (syndrom bits 1 5 7)
//  input bit  27 used 3 times (syndrom bits 3 5 6)
//  input bit  28 used 3 times (syndrom bits 1 3 4)
//  input bit  29 used 3 times (syndrom bits 0 2 5)
//  input bit  30 used 3 times (syndrom bits 0 3 8)
//  input bit  31 used 3 times (syndrom bits 1 2 8)
//  input bit  32 used 3 times (syndrom bits 2 4 6)
//  input bit  33 used 3 times (syndrom bits 4 7 8)
//  input bit  34 used 3 times (syndrom bits 1 6 7)
//  input bit  35 used 3 times (syndrom bits 0 3 5)
//  input bit  36 used 3 times (syndrom bits 0 3 7)
//  input bit  37 used 3 times (syndrom bits 1 5 6)
//  input bit  38 used 3 times (syndrom bits 2 4 8)
//  input bit  39 used 3 times (syndrom bits 1 4 8)
//  input bit  40 used 3 times (syndrom bits 2 5 6)
//  input bit  41 used 3 times (syndrom bits 0 3 6)
//  input bit  42 used 3 times (syndrom bits 0 5 7)
//  input bit  43 used 3 times (syndrom bits 2 3 7)
//  input bit  44 used 3 times (syndrom bits 3 4 8)
//  input bit  45 used 3 times (syndrom bits 1 4 7)
//  input bit  46 used 3 times (syndrom bits 1 7 8)
//  input bit  47 used 3 times (syndrom bits 0 2 6)
//  input bit  48 used 3 times (syndrom bits 2 5 8)
//  input bit  49 used 3 times (syndrom bits 0 5 6)
//  input bit  50 used 3 times (syndrom bits 1 4 5)
//  input bit  51 used 3 times (syndrom bits 0 1 3)
//  input bit  52 used 3 times (syndrom bits 2 3 4)
//  input bit  53 used 3 times (syndrom bits 3 6 8)
//  input bit  54 used 3 times (syndrom bits 0 6 7)
//  input bit  55 used 3 times (syndrom bits 2 7 8)
//  input bit  56 used 3 times (syndrom bits 1 2 4)
//  input bit  57 used 3 times (syndrom bits 4 5 7)
//  input bit  58 used 3 times (syndrom bits 0 1 5)
//  input bit  59 used 3 times (syndrom bits 5 6 8)
//  input bit  60 used 3 times (syndrom bits 1 3 8)
//  input bit  61 used 3 times (syndrom bits 2 3 6)
//  input bit  62 used 3 times (syndrom bits 0 4 6)
//  input bit  63 used 3 times (syndrom bits 0 7 8)
//  input bit  64 used 3 times (syndrom bits 3 4 7)
//  input bit  65 used 3 times (syndrom bits 1 2 7)
//  input bit  66 used 3 times (syndrom bits 2 4 5)
//  input bit  67 used 3 times (syndrom bits 3 5 8)
//  input bit  68 used 3 times (syndrom bits 0 1 6)
//  input bit  69 used 3 times (syndrom bits 0 1 4)
//  input bit  70 used 3 times (syndrom bits 5 6 7)
//  input bit  71 used 3 times (syndrom bits 2 3 8)
//  input bit  72 used 3 times (syndrom bits 3 7 8)
//  input bit  73 used 3 times (syndrom bits 2 6 8)
//  input bit  74 used 3 times (syndrom bits 0 4 5)
//  input bit  75 used 3 times (syndrom bits 0 1 7)
//  input bit  76 used 3 times (syndrom bits 1 4 6)
//  input bit  77 used 3 times (syndrom bits 2 3 5)
//  input bit  78 used 3 times (syndrom bits 4 5 6)
//  input bit  79 used 3 times (syndrom bits 1 2 3)
//  input bit  80 used 3 times (syndrom bits 0 5 8)
//  input bit  81 used 3 times (syndrom bits 2 4 7)
//  input bit  82 used 3 times (syndrom bits 1 3 7)
//  input bit  83 used 3 times (syndrom bits 0 6 8)
//  input bit  84 used 5 times (syndrom bits 0 3 6 7 8)
//  input bit  85 used 5 times (syndrom bits 0 1 2 4 5)
//  input bit  86 used 5 times (syndrom bits 1 2 4 5 8)
//  input bit  87 used 5 times (syndrom bits 1 2 3 6 7)
//  input bit  88 used 5 times (syndrom bits 3 4 5 6 7)
//  input bit  89 used 5 times (syndrom bits 0 4 6 7 8)
//  input bit  90 used 5 times (syndrom bits 0 1 3 5 8)
//  input bit  91 used 5 times (syndrom bits 0 2 3 5 8)
//  input bit  92 used 5 times (syndrom bits 1 2 4 6 7)
//  input bit  93 used 5 times (syndrom bits 1 2 6 7 8)
//  input bit  94 used 5 times (syndrom bits 0 2 3 4 5)
//  input bit  95 used 5 times (syndrom bits 0 1 3 4 5)
//  input bit  96 used 5 times (syndrom bits 3 4 6 7 8)
//  input bit  97 used 5 times (syndrom bits 0 5 6 7 8)
//  input bit  98 used 5 times (syndrom bits 0 1 2 6 7)
//  input bit  99 used 5 times (syndrom bits 1 2 3 5 8)
//  input bit 100 used 5 times (syndrom bits 1 2 3 4 8)
//  input bit 101 used 5 times (syndrom bits 0 4 5 6 7)
//  input bit 102 used 5 times (syndrom bits 1 4 5 6 7)
//  input bit 103 used 5 times (syndrom bits 0 2 3 4 8)
//  input bit 104 used 5 times (syndrom bits 0 2 3 6 8)
//  input bit 105 used 5 times (syndrom bits 0 1 2 5 7)
//  input bit 106 used 5 times (syndrom bits 1 3 5 7 8)
//  input bit 107 used 5 times (syndrom bits 4 5 6 7 8)
//  input bit 108 used 5 times (syndrom bits 0 1 3 4 6)
//  input bit 109 used 5 times (syndrom bits 1 2 3 4 6)
//  input bit 110 used 5 times (syndrom bits 0 2 5 7 8)
//  input bit 111 used 5 times (syndrom bits 0 2 5 6 7)
//  input bit 112 used 5 times (syndrom bits 0 1 3 4 8)
//  input bit 113 used 5 times (syndrom bits 1 3 4 5 8)
//  input bit 114 used 5 times (syndrom bits 2 4 6 7 8)
//  input bit 115 used 5 times (syndrom bits 1 2 5 6 7)
//  input bit 116 used 5 times (syndrom bits 0 2 3 6 7)
//  input bit 117 used 5 times (syndrom bits 0 1 2 3 5)
//  input bit 118 used 5 times (syndrom bits 0 3 4 5 8)
//  input bit 119 used 5 times (syndrom bits 1 4 6 7 8)
//  input bit 120 used 5 times (syndrom bits 1 3 4 7 8)
//  input bit 121 used 5 times (syndrom bits 0 2 5 6 8)
//  input bit 122 used 5 times (syndrom bits 0 2 4 5 6)
//  input bit 123 used 5 times (syndrom bits 0 1 3 6 7)
//  input bit 124 used 5 times (syndrom bits 1 2 3 5 7)
//  input bit 125 used 5 times (syndrom bits 1 4 5 7 8)
//  input bit 126 used 5 times (syndrom bits 2 3 4 6 8)
//  input bit 127 used 5 times (syndrom bits 0 3 4 6 8)
function [9-1:0] extended_hamming_code_137_128_f;
    input [128-1:0] in;
    reg [9-1:0] syndrom;
    begin
        syndrom[0] = in[  0]^in[  5]^in[  6]^in[ 11]^in[ 12]^in[ 17]^in[ 18]^in[ 23]^in[ 24]^in[ 29]^in[ 30]^in[ 35]^in[ 36]^in[ 41]^in[ 42]^in[ 47]^in[ 49]^in[ 51]^in[ 54]^in[ 58]^in[ 62]^in[ 63]^in[ 68]^in[ 69]^in[ 74]^in[ 75]^in[ 80]^in[ 83]^in[ 84]^in[ 85]^in[ 89]^in[ 90]^in[ 91]^in[ 94]^in[ 95]^in[ 97]^in[ 98]^in[101]^in[103]^in[104]^in[105]^in[108]^in[110]^in[111]^in[112]^in[116]^in[117]^in[118]^in[121]^in[122]^in[123]^in[127];//52 inputs
        syndrom[1] = in[  0]^in[  5]^in[  7]^in[  9]^in[ 14]^in[ 15]^in[ 20]^in[ 21]^in[ 26]^in[ 28]^in[ 31]^in[ 34]^in[ 37]^in[ 39]^in[ 45]^in[ 46]^in[ 50]^in[ 51]^in[ 56]^in[ 58]^in[ 60]^in[ 65]^in[ 68]^in[ 69]^in[ 75]^in[ 76]^in[ 79]^in[ 82]^in[ 85]^in[ 86]^in[ 87]^in[ 90]^in[ 92]^in[ 93]^in[ 95]^in[ 98]^in[ 99]^in[100]^in[102]^in[105]^in[106]^in[108]^in[109]^in[112]^in[113]^in[115]^in[117]^in[119]^in[120]^in[123]^in[124]^in[125];//52 inputs
        syndrom[2] = in[  0]^in[  6]^in[  7]^in[  8]^in[ 14]^in[ 16]^in[ 18]^in[ 23]^in[ 24]^in[ 29]^in[ 31]^in[ 32]^in[ 38]^in[ 40]^in[ 43]^in[ 47]^in[ 48]^in[ 52]^in[ 55]^in[ 56]^in[ 61]^in[ 65]^in[ 66]^in[ 71]^in[ 73]^in[ 77]^in[ 79]^in[ 81]^in[ 85]^in[ 86]^in[ 87]^in[ 91]^in[ 92]^in[ 93]^in[ 94]^in[ 98]^in[ 99]^in[100]^in[103]^in[104]^in[105]^in[109]^in[110]^in[111]^in[114]^in[115]^in[116]^in[117]^in[121]^in[122]^in[124]^in[126];//52 inputs
        syndrom[3] = in[  1]^in[  3]^in[  9]^in[ 10]^in[ 12]^in[ 18]^in[ 19]^in[ 21]^in[ 27]^in[ 28]^in[ 30]^in[ 35]^in[ 36]^in[ 41]^in[ 43]^in[ 44]^in[ 51]^in[ 52]^in[ 53]^in[ 60]^in[ 61]^in[ 64]^in[ 67]^in[ 71]^in[ 72]^in[ 77]^in[ 79]^in[ 82]^in[ 84]^in[ 87]^in[ 88]^in[ 90]^in[ 91]^in[ 94]^in[ 95]^in[ 96]^in[ 99]^in[100]^in[103]^in[104]^in[106]^in[108]^in[109]^in[112]^in[113]^in[116]^in[117]^in[118]^in[120]^in[123]^in[124]^in[126]^in[127];//53 inputs
        syndrom[4] = in[  1]^in[  4]^in[  6]^in[ 11]^in[ 12]^in[ 17]^in[ 19]^in[ 22]^in[ 25]^in[ 28]^in[ 32]^in[ 33]^in[ 38]^in[ 39]^in[ 44]^in[ 45]^in[ 50]^in[ 52]^in[ 56]^in[ 57]^in[ 62]^in[ 64]^in[ 66]^in[ 69]^in[ 74]^in[ 76]^in[ 78]^in[ 81]^in[ 85]^in[ 86]^in[ 88]^in[ 89]^in[ 92]^in[ 94]^in[ 95]^in[ 96]^in[100]^in[101]^in[102]^in[103]^in[107]^in[108]^in[109]^in[112]^in[113]^in[114]^in[118]^in[119]^in[120]^in[122]^in[125]^in[126]^in[127];//53 inputs
        syndrom[5] = in[  1]^in[  4]^in[  7]^in[ 10]^in[ 13]^in[ 16]^in[ 20]^in[ 21]^in[ 26]^in[ 27]^in[ 29]^in[ 35]^in[ 37]^in[ 40]^in[ 42]^in[ 48]^in[ 49]^in[ 50]^in[ 57]^in[ 58]^in[ 59]^in[ 66]^in[ 67]^in[ 70]^in[ 74]^in[ 77]^in[ 78]^in[ 80]^in[ 85]^in[ 86]^in[ 88]^in[ 90]^in[ 91]^in[ 94]^in[ 95]^in[ 97]^in[ 99]^in[101]^in[102]^in[105]^in[106]^in[107]^in[110]^in[111]^in[113]^in[115]^in[117]^in[118]^in[121]^in[122]^in[124]^in[125];//52 inputs
        syndrom[6] = in[  2]^in[  3]^in[  8]^in[  9]^in[ 14]^in[ 15]^in[ 19]^in[ 22]^in[ 25]^in[ 27]^in[ 32]^in[ 34]^in[ 37]^in[ 40]^in[ 41]^in[ 47]^in[ 49]^in[ 53]^in[ 54]^in[ 59]^in[ 61]^in[ 62]^in[ 68]^in[ 70]^in[ 73]^in[ 76]^in[ 78]^in[ 83]^in[ 84]^in[ 87]^in[ 88]^in[ 89]^in[ 92]^in[ 93]^in[ 96]^in[ 97]^in[ 98]^in[101]^in[102]^in[104]^in[107]^in[108]^in[109]^in[111]^in[114]^in[115]^in[116]^in[119]^in[121]^in[122]^in[123]^in[126]^in[127];//53 inputs
        syndrom[7] = in[  2]^in[  3]^in[  8]^in[ 10]^in[ 13]^in[ 16]^in[ 17]^in[ 23]^in[ 25]^in[ 26]^in[ 33]^in[ 34]^in[ 36]^in[ 42]^in[ 43]^in[ 45]^in[ 46]^in[ 54]^in[ 55]^in[ 57]^in[ 63]^in[ 64]^in[ 65]^in[ 70]^in[ 72]^in[ 75]^in[ 81]^in[ 82]^in[ 84]^in[ 87]^in[ 88]^in[ 89]^in[ 92]^in[ 93]^in[ 96]^in[ 97]^in[ 98]^in[101]^in[102]^in[105]^in[106]^in[107]^in[110]^in[111]^in[114]^in[115]^in[116]^in[119]^in[120]^in[123]^in[124]^in[125];//52 inputs
        syndrom[8] = in[  2]^in[  4]^in[  5]^in[ 11]^in[ 13]^in[ 15]^in[ 20]^in[ 22]^in[ 24]^in[ 30]^in[ 31]^in[ 33]^in[ 38]^in[ 39]^in[ 44]^in[ 46]^in[ 48]^in[ 53]^in[ 55]^in[ 59]^in[ 60]^in[ 63]^in[ 67]^in[ 71]^in[ 72]^in[ 73]^in[ 80]^in[ 83]^in[ 84]^in[ 86]^in[ 89]^in[ 90]^in[ 91]^in[ 93]^in[ 96]^in[ 97]^in[ 99]^in[100]^in[103]^in[104]^in[106]^in[107]^in[110]^in[112]^in[113]^in[114]^in[118]^in[119]^in[120]^in[121]^in[125]^in[126]^in[127];//53 inputs
        extended_hamming_code_137_128_f = syndrom;
    end
endfunction
function [2+128-1:0] extended_hamming_code_137_128_f_correction_pattern_f;
    input [9-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [128-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {128{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			9'b000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {128{1'b0}};
			end	
			9'b000000111: begin
				correction_pattern = {128{1'b0}};correction_pattern[  0]=1'b1;
			end
			9'b000111000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  1]=1'b1;
			end
			9'b111000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  2]=1'b1;
			end
			9'b011001000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  3]=1'b1;
			end
			9'b100110000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  4]=1'b1;
			end
			9'b100000011: begin
				correction_pattern = {128{1'b0}};correction_pattern[  5]=1'b1;
			end
			9'b000010101: begin
				correction_pattern = {128{1'b0}};correction_pattern[  6]=1'b1;
			end
			9'b000100110: begin
				correction_pattern = {128{1'b0}};correction_pattern[  7]=1'b1;
			end
			9'b011000100: begin
				correction_pattern = {128{1'b0}};correction_pattern[  8]=1'b1;
			end
			9'b001001010: begin
				correction_pattern = {128{1'b0}};correction_pattern[  9]=1'b1;
			end
			9'b010101000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 10]=1'b1;
			end
			9'b100010001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 11]=1'b1;
			end
			9'b000011001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 12]=1'b1;
			end
			9'b110100000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 13]=1'b1;
			end
			9'b001000110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 14]=1'b1;
			end
			9'b101000010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 15]=1'b1;
			end
			9'b010100100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 16]=1'b1;
			end
			9'b010010001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 17]=1'b1;
			end
			9'b000001101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 18]=1'b1;
			end
			9'b001011000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 19]=1'b1;
			end
			9'b100100010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 20]=1'b1;
			end
			9'b000101010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 21]=1'b1;
			end
			9'b101010000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 22]=1'b1;
			end
			9'b010000101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 23]=1'b1;
			end
			9'b100000101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 24]=1'b1;
			end
			9'b011010000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 25]=1'b1;
			end
			9'b010100010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 26]=1'b1;
			end
			9'b001101000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 27]=1'b1;
			end
			9'b000011010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 28]=1'b1;
			end
			9'b000100101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 29]=1'b1;
			end
			9'b100001001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 30]=1'b1;
			end
			9'b100000110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 31]=1'b1;
			end
			9'b001010100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 32]=1'b1;
			end
			9'b110010000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 33]=1'b1;
			end
			9'b011000010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 34]=1'b1;
			end
			9'b000101001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 35]=1'b1;
			end
			9'b010001001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 36]=1'b1;
			end
			9'b001100010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 37]=1'b1;
			end
			9'b100010100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 38]=1'b1;
			end
			9'b100010010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 39]=1'b1;
			end
			9'b001100100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 40]=1'b1;
			end
			9'b001001001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 41]=1'b1;
			end
			9'b010100001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 42]=1'b1;
			end
			9'b010001100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 43]=1'b1;
			end
			9'b100011000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 44]=1'b1;
			end
			9'b010010010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 45]=1'b1;
			end
			9'b110000010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 46]=1'b1;
			end
			9'b001000101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 47]=1'b1;
			end
			9'b100100100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 48]=1'b1;
			end
			9'b001100001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 49]=1'b1;
			end
			9'b000110010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 50]=1'b1;
			end
			9'b000001011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 51]=1'b1;
			end
			9'b000011100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 52]=1'b1;
			end
			9'b101001000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 53]=1'b1;
			end
			9'b011000001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 54]=1'b1;
			end
			9'b110000100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 55]=1'b1;
			end
			9'b000010110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 56]=1'b1;
			end
			9'b010110000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 57]=1'b1;
			end
			9'b000100011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 58]=1'b1;
			end
			9'b101100000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 59]=1'b1;
			end
			9'b100001010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 60]=1'b1;
			end
			9'b001001100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 61]=1'b1;
			end
			9'b001010001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 62]=1'b1;
			end
			9'b110000001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 63]=1'b1;
			end
			9'b010011000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 64]=1'b1;
			end
			9'b010000110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 65]=1'b1;
			end
			9'b000110100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 66]=1'b1;
			end
			9'b100101000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 67]=1'b1;
			end
			9'b001000011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 68]=1'b1;
			end
			9'b000010011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 69]=1'b1;
			end
			9'b011100000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 70]=1'b1;
			end
			9'b100001100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 71]=1'b1;
			end
			9'b110001000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 72]=1'b1;
			end
			9'b101000100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 73]=1'b1;
			end
			9'b000110001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 74]=1'b1;
			end
			9'b010000011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 75]=1'b1;
			end
			9'b001010010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 76]=1'b1;
			end
			9'b000101100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 77]=1'b1;
			end
			9'b001110000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 78]=1'b1;
			end
			9'b000001110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 79]=1'b1;
			end
			9'b100100001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 80]=1'b1;
			end
			9'b010010100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 81]=1'b1;
			end
			9'b010001010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 82]=1'b1;
			end
			9'b101000001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 83]=1'b1;
			end
			9'b111001001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 84]=1'b1;
			end
			9'b000110111: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 85]=1'b1;
			end
			9'b100110110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 86]=1'b1;
			end
			9'b011001110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 87]=1'b1;
			end
			9'b011111000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 88]=1'b1;
			end
			9'b111010001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 89]=1'b1;
			end
			9'b100101011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 90]=1'b1;
			end
			9'b100101101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 91]=1'b1;
			end
			9'b011010110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 92]=1'b1;
			end
			9'b111000110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 93]=1'b1;
			end
			9'b000111101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 94]=1'b1;
			end
			9'b000111011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 95]=1'b1;
			end
			9'b111011000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 96]=1'b1;
			end
			9'b111100001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 97]=1'b1;
			end
			9'b011000111: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 98]=1'b1;
			end
			9'b100101110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 99]=1'b1;
			end
			9'b100011110: begin
				correction_pattern = {128{1'b0}};correction_pattern[100]=1'b1;
			end
			9'b011110001: begin
				correction_pattern = {128{1'b0}};correction_pattern[101]=1'b1;
			end
			9'b011110010: begin
				correction_pattern = {128{1'b0}};correction_pattern[102]=1'b1;
			end
			9'b100011101: begin
				correction_pattern = {128{1'b0}};correction_pattern[103]=1'b1;
			end
			9'b101001101: begin
				correction_pattern = {128{1'b0}};correction_pattern[104]=1'b1;
			end
			9'b010100111: begin
				correction_pattern = {128{1'b0}};correction_pattern[105]=1'b1;
			end
			9'b110101010: begin
				correction_pattern = {128{1'b0}};correction_pattern[106]=1'b1;
			end
			9'b111110000: begin
				correction_pattern = {128{1'b0}};correction_pattern[107]=1'b1;
			end
			9'b001011011: begin
				correction_pattern = {128{1'b0}};correction_pattern[108]=1'b1;
			end
			9'b001011110: begin
				correction_pattern = {128{1'b0}};correction_pattern[109]=1'b1;
			end
			9'b110100101: begin
				correction_pattern = {128{1'b0}};correction_pattern[110]=1'b1;
			end
			9'b011100101: begin
				correction_pattern = {128{1'b0}};correction_pattern[111]=1'b1;
			end
			9'b100011011: begin
				correction_pattern = {128{1'b0}};correction_pattern[112]=1'b1;
			end
			9'b100111010: begin
				correction_pattern = {128{1'b0}};correction_pattern[113]=1'b1;
			end
			9'b111010100: begin
				correction_pattern = {128{1'b0}};correction_pattern[114]=1'b1;
			end
			9'b011100110: begin
				correction_pattern = {128{1'b0}};correction_pattern[115]=1'b1;
			end
			9'b011001101: begin
				correction_pattern = {128{1'b0}};correction_pattern[116]=1'b1;
			end
			9'b000101111: begin
				correction_pattern = {128{1'b0}};correction_pattern[117]=1'b1;
			end
			9'b100111001: begin
				correction_pattern = {128{1'b0}};correction_pattern[118]=1'b1;
			end
			9'b111010010: begin
				correction_pattern = {128{1'b0}};correction_pattern[119]=1'b1;
			end
			9'b110011010: begin
				correction_pattern = {128{1'b0}};correction_pattern[120]=1'b1;
			end
			9'b101100101: begin
				correction_pattern = {128{1'b0}};correction_pattern[121]=1'b1;
			end
			9'b001110101: begin
				correction_pattern = {128{1'b0}};correction_pattern[122]=1'b1;
			end
			9'b011001011: begin
				correction_pattern = {128{1'b0}};correction_pattern[123]=1'b1;
			end
			9'b010101110: begin
				correction_pattern = {128{1'b0}};correction_pattern[124]=1'b1;
			end
			9'b110110010: begin
				correction_pattern = {128{1'b0}};correction_pattern[125]=1'b1;
			end
			9'b101011100: begin
				correction_pattern = {128{1'b0}};correction_pattern[126]=1'b1;
			end
			9'b101011001: begin
				correction_pattern = {128{1'b0}};correction_pattern[127]=1'b1;
			end
			9'b000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			9'b100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_137_128_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [9-1:0] stored_data_edc = extended_hamming_code_137_128_f(i_stored_data);
wire [9-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [128-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_137_128_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule


/////////////////////////////////////////////////////////////////////////////////////////////////
// *_min_delay modules: use the least logic gates between input and outputs (keep logic shallow)
/////////////////////////////////////////////////////////////////////////////////////////////////
module edc_hc_4_min_delay (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: x x  (2 inputs)
//  syndrom[1]: x  x (2 inputs)
//  syndrom[2]:  xx  (2 inputs)
//  syndrom[3]:  x x (2 inputs)
//Input usage report:
//  input bit 0 used 2 times (syndrom bits 0 1)
//  input bit 1 used 2 times (syndrom bits 2 3)
//  input bit 2 used 2 times (syndrom bits 0 2)
//  input bit 3 used 2 times (syndrom bits 1 3)
function [4-1:0] hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[2];//2 inputs
        syndrom[1] = in[0]^in[3];//2 inputs
        syndrom[2] = in[1]^in[2];//2 inputs
        syndrom[3] = in[1]^in[3];//2 inputs
        hamming_code_8_4_f = syndrom;
    end
endfunction
wire [4-1:0] stored_data_edc = hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_4_min_delay (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: xxx  (3 inputs)
//  syndrom[1]: xx x (3 inputs)
//  syndrom[2]: x xx (3 inputs)
//  syndrom[3]:  xxx (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 1 3)
//  input bit 2 used 3 times (syndrom bits 0 2 3)
//  input bit 3 used 3 times (syndrom bits 1 2 3)
function [4-1:0] extended_hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[2];//3 inputs
        syndrom[1] = in[0]^in[1]^in[3];//3 inputs
        syndrom[2] = in[0]^in[2]^in[3];//3 inputs
        syndrom[3] = in[1]^in[2]^in[3];//3 inputs
        extended_hamming_code_8_4_f = syndrom;
    end
endfunction
wire [4-1:0] stored_data_edc = extended_hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_4_min_delay (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [4-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: xxx  (3 inputs)
//  syndrom[1]: xx x (3 inputs)
//  syndrom[2]: x xx (3 inputs)
//  syndrom[3]:  xxx (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 1 3)
//  input bit 2 used 3 times (syndrom bits 0 2 3)
//  input bit 3 used 3 times (syndrom bits 1 2 3)
function [4-1:0] extended_hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[2];//3 inputs
        syndrom[1] = in[0]^in[1]^in[3];//3 inputs
        syndrom[2] = in[0]^in[2]^in[3];//3 inputs
        syndrom[3] = in[1]^in[2]^in[3];//3 inputs
        extended_hamming_code_8_4_f = syndrom;
    end
endfunction
function [2+4-1:0] extended_hamming_code_8_4_f_correction_pattern_f;
    input [4-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [4-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {4{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			4'b0000: begin
				correctable_error = 1'b0;
				correction_pattern = {4{1'b0}};
			end	
			4'b0111: begin
				correction_pattern = {4{1'b0}};correction_pattern[0]=1'b1;
			end
			4'b1011: begin
				correction_pattern = {4{1'b0}};correction_pattern[1]=1'b1;
			end
			4'b1101: begin
				correction_pattern = {4{1'b0}};correction_pattern[2]=1'b1;
			end
			4'b1110: begin
				correction_pattern = {4{1'b0}};correction_pattern[3]=1'b1;
			end
			4'b0001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b0010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b0100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b1000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_8_4_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [4-1:0] stored_data_edc = extended_hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [4-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_8_4_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_8_min_delay (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_16_8_f
//Compute 8 bits Error Detection Code from a 8 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 256 valid code words out of 65536 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: x     x  (2 inputs)
//  syndrom[1]: x      x (2 inputs)
//  syndrom[2]:  x    x  (2 inputs)
//  syndrom[3]:  x     x (2 inputs)
//  syndrom[4]:   x x    (2 inputs)
//  syndrom[5]:   x  x   (2 inputs)
//  syndrom[6]:    xx    (2 inputs)
//  syndrom[7]:    x x   (2 inputs)
//Input usage report:
//  input bit 0 used 2 times (syndrom bits 0 1)
//  input bit 1 used 2 times (syndrom bits 2 3)
//  input bit 2 used 2 times (syndrom bits 4 5)
//  input bit 3 used 2 times (syndrom bits 6 7)
//  input bit 4 used 2 times (syndrom bits 4 6)
//  input bit 5 used 2 times (syndrom bits 5 7)
//  input bit 6 used 2 times (syndrom bits 0 2)
//  input bit 7 used 2 times (syndrom bits 1 3)
function [8-1:0] hamming_code_16_8_f;
    input [8-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[6];//2 inputs
        syndrom[1] = in[0]^in[7];//2 inputs
        syndrom[2] = in[1]^in[6];//2 inputs
        syndrom[3] = in[1]^in[7];//2 inputs
        syndrom[4] = in[2]^in[4];//2 inputs
        syndrom[5] = in[2]^in[5];//2 inputs
        syndrom[6] = in[3]^in[4];//2 inputs
        syndrom[7] = in[3]^in[5];//2 inputs
        hamming_code_16_8_f = syndrom;
    end
endfunction
wire [8-1:0] stored_data_edc = hamming_code_16_8_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_8_min_delay (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_16_8_f
//Compute 8 bits Error Detection Code from a 8 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 256 valid code words out of 65536 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: x   xx   (3 inputs)
//  syndrom[1]: x   x x  (3 inputs)
//  syndrom[2]: x    xx  (3 inputs)
//  syndrom[3]:  xx    x (3 inputs)
//  syndrom[4]:  x x   x (3 inputs)
//  syndrom[5]:  x  xx   (3 inputs)
//  syndrom[6]:   xx  x  (3 inputs)
//  syndrom[7]:   xx   x (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 3 4 5)
//  input bit 2 used 3 times (syndrom bits 3 6 7)
//  input bit 3 used 3 times (syndrom bits 4 6 7)
//  input bit 4 used 3 times (syndrom bits 0 1 5)
//  input bit 5 used 3 times (syndrom bits 0 2 5)
//  input bit 6 used 3 times (syndrom bits 1 2 6)
//  input bit 7 used 3 times (syndrom bits 3 4 7)
function [8-1:0] extended_hamming_code_16_8_f;
    input [8-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[4]^in[5];//3 inputs
        syndrom[1] = in[0]^in[4]^in[6];//3 inputs
        syndrom[2] = in[0]^in[5]^in[6];//3 inputs
        syndrom[3] = in[1]^in[2]^in[7];//3 inputs
        syndrom[4] = in[1]^in[3]^in[7];//3 inputs
        syndrom[5] = in[1]^in[4]^in[5];//3 inputs
        syndrom[6] = in[2]^in[3]^in[6];//3 inputs
        syndrom[7] = in[2]^in[3]^in[7];//3 inputs
        extended_hamming_code_16_8_f = syndrom;
    end
endfunction
wire [8-1:0] stored_data_edc = extended_hamming_code_16_8_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_8_min_delay (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [8-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_16_8_f
//Compute 8 bits Error Detection Code from a 8 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 256 valid code words out of 65536 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: x   xx   (3 inputs)
//  syndrom[1]: x   x x  (3 inputs)
//  syndrom[2]: x    xx  (3 inputs)
//  syndrom[3]:  xx    x (3 inputs)
//  syndrom[4]:  x x   x (3 inputs)
//  syndrom[5]:  x  xx   (3 inputs)
//  syndrom[6]:   xx  x  (3 inputs)
//  syndrom[7]:   xx   x (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 3 4 5)
//  input bit 2 used 3 times (syndrom bits 3 6 7)
//  input bit 3 used 3 times (syndrom bits 4 6 7)
//  input bit 4 used 3 times (syndrom bits 0 1 5)
//  input bit 5 used 3 times (syndrom bits 0 2 5)
//  input bit 6 used 3 times (syndrom bits 1 2 6)
//  input bit 7 used 3 times (syndrom bits 3 4 7)
function [8-1:0] extended_hamming_code_16_8_f;
    input [8-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[4]^in[5];//3 inputs
        syndrom[1] = in[0]^in[4]^in[6];//3 inputs
        syndrom[2] = in[0]^in[5]^in[6];//3 inputs
        syndrom[3] = in[1]^in[2]^in[7];//3 inputs
        syndrom[4] = in[1]^in[3]^in[7];//3 inputs
        syndrom[5] = in[1]^in[4]^in[5];//3 inputs
        syndrom[6] = in[2]^in[3]^in[6];//3 inputs
        syndrom[7] = in[2]^in[3]^in[7];//3 inputs
        extended_hamming_code_16_8_f = syndrom;
    end
endfunction
function [2+8-1:0] extended_hamming_code_16_8_f_correction_pattern_f;
    input [8-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [8-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {8{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			8'b00000000: begin
				correctable_error = 1'b0;
				correction_pattern = {8{1'b0}};
			end	
			8'b00000111: begin
				correction_pattern = {8{1'b0}};correction_pattern[0]=1'b1;
			end
			8'b00111000: begin
				correction_pattern = {8{1'b0}};correction_pattern[1]=1'b1;
			end
			8'b11001000: begin
				correction_pattern = {8{1'b0}};correction_pattern[2]=1'b1;
			end
			8'b11010000: begin
				correction_pattern = {8{1'b0}};correction_pattern[3]=1'b1;
			end
			8'b00100011: begin
				correction_pattern = {8{1'b0}};correction_pattern[4]=1'b1;
			end
			8'b00100101: begin
				correction_pattern = {8{1'b0}};correction_pattern[5]=1'b1;
			end
			8'b01000110: begin
				correction_pattern = {8{1'b0}};correction_pattern[6]=1'b1;
			end
			8'b10011000: begin
				correction_pattern = {8{1'b0}};correction_pattern[7]=1'b1;
			end
			8'b00000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b01000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b10000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_16_8_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [8-1:0] stored_data_edc = extended_hamming_code_16_8_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [8-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_16_8_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_12_min_delay (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [12-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [12-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_24_12_f
//Compute 12 bits Error Detection Code from a 12 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 16777216 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[ 0]: x         x  (2 inputs)
//  syndrom[ 1]: x          x (2 inputs)
//  syndrom[ 2]:  x        x  (2 inputs)
//  syndrom[ 3]:  x         x (2 inputs)
//  syndrom[ 4]:   x     x    (2 inputs)
//  syndrom[ 5]:   x      x   (2 inputs)
//  syndrom[ 6]:    x    x    (2 inputs)
//  syndrom[ 7]:    x     x   (2 inputs)
//  syndrom[ 8]:     x x      (2 inputs)
//  syndrom[ 9]:     x  x     (2 inputs)
//  syndrom[10]:      xx      (2 inputs)
//  syndrom[11]:      x x     (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 8 10)
//  input bit  7 used  2 times (syndrom bits 9 11)
//  input bit  8 used  2 times (syndrom bits 4 6)
//  input bit  9 used  2 times (syndrom bits 5 7)
//  input bit 10 used  2 times (syndrom bits 0 2)
//  input bit 11 used  2 times (syndrom bits 1 3)
function [12-1:0] hamming_code_24_12_f;
    input [12-1:0] in;
    reg [12-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[10];//2 inputs
        syndrom[ 1] = in[ 0]^in[11];//2 inputs
        syndrom[ 2] = in[ 1]^in[10];//2 inputs
        syndrom[ 3] = in[ 1]^in[11];//2 inputs
        syndrom[ 4] = in[ 2]^in[ 8];//2 inputs
        syndrom[ 5] = in[ 2]^in[ 9];//2 inputs
        syndrom[ 6] = in[ 3]^in[ 8];//2 inputs
        syndrom[ 7] = in[ 3]^in[ 9];//2 inputs
        syndrom[ 8] = in[ 4]^in[ 6];//2 inputs
        syndrom[ 9] = in[ 4]^in[ 7];//2 inputs
        syndrom[10] = in[ 5]^in[ 6];//2 inputs
        syndrom[11] = in[ 5]^in[ 7];//2 inputs
        hamming_code_24_12_f = syndrom;
    end
endfunction
wire [12-1:0] stored_data_edc = hamming_code_24_12_f(i_stored_data);
wire [12-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_12_min_delay (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [12-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [12-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_24_12_f
//Compute 12 bits Error Detection Code from a 12 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 16777216 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[ 0]: x     x  x   (3 inputs)
//  syndrom[ 1]: x      xx    (3 inputs)
//  syndrom[ 2]: x      x x   (3 inputs)
//  syndrom[ 3]:  x    x x    (3 inputs)
//  syndrom[ 4]:  x    x  x   (3 inputs)
//  syndrom[ 5]:  x     xx    (3 inputs)
//  syndrom[ 6]:   x x      x (3 inputs)
//  syndrom[ 7]:   x  x    x  (3 inputs)
//  syndrom[ 8]:   x  x     x (3 inputs)
//  syndrom[ 9]:    xx     x  (3 inputs)
//  syndrom[10]:    xx      x (3 inputs)
//  syndrom[11]:    x x    x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 6 9 10)
//  input bit  5 used  3 times (syndrom bits 7 8 11)
//  input bit  6 used  3 times (syndrom bits 0 3 4)
//  input bit  7 used  3 times (syndrom bits 1 2 5)
//  input bit  8 used  3 times (syndrom bits 1 3 5)
//  input bit  9 used  3 times (syndrom bits 0 2 4)
//  input bit 10 used  3 times (syndrom bits 7 9 11)
//  input bit 11 used  3 times (syndrom bits 6 8 10)
function [12-1:0] extended_hamming_code_24_12_f;
    input [12-1:0] in;
    reg [12-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 6]^in[ 9];//3 inputs
        syndrom[ 1] = in[ 0]^in[ 7]^in[ 8];//3 inputs
        syndrom[ 2] = in[ 0]^in[ 7]^in[ 9];//3 inputs
        syndrom[ 3] = in[ 1]^in[ 6]^in[ 8];//3 inputs
        syndrom[ 4] = in[ 1]^in[ 6]^in[ 9];//3 inputs
        syndrom[ 5] = in[ 1]^in[ 7]^in[ 8];//3 inputs
        syndrom[ 6] = in[ 2]^in[ 4]^in[11];//3 inputs
        syndrom[ 7] = in[ 2]^in[ 5]^in[10];//3 inputs
        syndrom[ 8] = in[ 2]^in[ 5]^in[11];//3 inputs
        syndrom[ 9] = in[ 3]^in[ 4]^in[10];//3 inputs
        syndrom[10] = in[ 3]^in[ 4]^in[11];//3 inputs
        syndrom[11] = in[ 3]^in[ 5]^in[10];//3 inputs
        extended_hamming_code_24_12_f = syndrom;
    end
endfunction
wire [12-1:0] stored_data_edc = extended_hamming_code_24_12_f(i_stored_data);
wire [12-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_12_min_delay (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [12-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [12-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [12-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_24_12_f
//Compute 12 bits Error Detection Code from a 12 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 16777216 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[ 0]: x     x  x   (3 inputs)
//  syndrom[ 1]: x      xx    (3 inputs)
//  syndrom[ 2]: x      x x   (3 inputs)
//  syndrom[ 3]:  x    x x    (3 inputs)
//  syndrom[ 4]:  x    x  x   (3 inputs)
//  syndrom[ 5]:  x     xx    (3 inputs)
//  syndrom[ 6]:   x x      x (3 inputs)
//  syndrom[ 7]:   x  x    x  (3 inputs)
//  syndrom[ 8]:   x  x     x (3 inputs)
//  syndrom[ 9]:    xx     x  (3 inputs)
//  syndrom[10]:    xx      x (3 inputs)
//  syndrom[11]:    x x    x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 6 9 10)
//  input bit  5 used  3 times (syndrom bits 7 8 11)
//  input bit  6 used  3 times (syndrom bits 0 3 4)
//  input bit  7 used  3 times (syndrom bits 1 2 5)
//  input bit  8 used  3 times (syndrom bits 1 3 5)
//  input bit  9 used  3 times (syndrom bits 0 2 4)
//  input bit 10 used  3 times (syndrom bits 7 9 11)
//  input bit 11 used  3 times (syndrom bits 6 8 10)
function [12-1:0] extended_hamming_code_24_12_f;
    input [12-1:0] in;
    reg [12-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 6]^in[ 9];//3 inputs
        syndrom[ 1] = in[ 0]^in[ 7]^in[ 8];//3 inputs
        syndrom[ 2] = in[ 0]^in[ 7]^in[ 9];//3 inputs
        syndrom[ 3] = in[ 1]^in[ 6]^in[ 8];//3 inputs
        syndrom[ 4] = in[ 1]^in[ 6]^in[ 9];//3 inputs
        syndrom[ 5] = in[ 1]^in[ 7]^in[ 8];//3 inputs
        syndrom[ 6] = in[ 2]^in[ 4]^in[11];//3 inputs
        syndrom[ 7] = in[ 2]^in[ 5]^in[10];//3 inputs
        syndrom[ 8] = in[ 2]^in[ 5]^in[11];//3 inputs
        syndrom[ 9] = in[ 3]^in[ 4]^in[10];//3 inputs
        syndrom[10] = in[ 3]^in[ 4]^in[11];//3 inputs
        syndrom[11] = in[ 3]^in[ 5]^in[10];//3 inputs
        extended_hamming_code_24_12_f = syndrom;
    end
endfunction
function [2+12-1:0] extended_hamming_code_24_12_f_correction_pattern_f;
    input [12-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [12-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {12{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			12'b000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {12{1'b0}};
			end	
			12'b000000000111: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 0]=1'b1;
			end
			12'b000000111000: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 1]=1'b1;
			end
			12'b000111000000: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 2]=1'b1;
			end
			12'b111000000000: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 3]=1'b1;
			end
			12'b011001000000: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 4]=1'b1;
			end
			12'b100110000000: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 5]=1'b1;
			end
			12'b000000011001: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 6]=1'b1;
			end
			12'b000000100110: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 7]=1'b1;
			end
			12'b000000101010: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 8]=1'b1;
			end
			12'b000000010101: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 9]=1'b1;
			end
			12'b101010000000: begin
				correction_pattern = {12{1'b0}};correction_pattern[10]=1'b1;
			end
			12'b010101000000: begin
				correction_pattern = {12{1'b0}};correction_pattern[11]=1'b1;
			end
			12'b000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_24_12_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [12-1:0] stored_data_edc = extended_hamming_code_24_12_f(i_stored_data);
wire [12-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [12-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_24_12_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_16_min_delay (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [16-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [16-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_32_16_f
//Compute 16 bits Error Detection Code from a 16 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 4294967296 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[ 0]: x             x  (2 inputs)
//  syndrom[ 1]: x              x (2 inputs)
//  syndrom[ 2]:  x            x  (2 inputs)
//  syndrom[ 3]:  x             x (2 inputs)
//  syndrom[ 4]:   x         x    (2 inputs)
//  syndrom[ 5]:   x          x   (2 inputs)
//  syndrom[ 6]:    x        x    (2 inputs)
//  syndrom[ 7]:    x         x   (2 inputs)
//  syndrom[ 8]:     x     x      (2 inputs)
//  syndrom[ 9]:     x      x     (2 inputs)
//  syndrom[10]:      x    x      (2 inputs)
//  syndrom[11]:      x     x     (2 inputs)
//  syndrom[12]:       x x        (2 inputs)
//  syndrom[13]:       x  x       (2 inputs)
//  syndrom[14]:        xx        (2 inputs)
//  syndrom[15]:        x x       (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 12 14)
//  input bit  9 used  2 times (syndrom bits 13 15)
//  input bit 10 used  2 times (syndrom bits 8 10)
//  input bit 11 used  2 times (syndrom bits 9 11)
//  input bit 12 used  2 times (syndrom bits 4 6)
//  input bit 13 used  2 times (syndrom bits 5 7)
//  input bit 14 used  2 times (syndrom bits 0 2)
//  input bit 15 used  2 times (syndrom bits 1 3)
function [16-1:0] hamming_code_32_16_f;
    input [16-1:0] in;
    reg [16-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[14];//2 inputs
        syndrom[ 1] = in[ 0]^in[15];//2 inputs
        syndrom[ 2] = in[ 1]^in[14];//2 inputs
        syndrom[ 3] = in[ 1]^in[15];//2 inputs
        syndrom[ 4] = in[ 2]^in[12];//2 inputs
        syndrom[ 5] = in[ 2]^in[13];//2 inputs
        syndrom[ 6] = in[ 3]^in[12];//2 inputs
        syndrom[ 7] = in[ 3]^in[13];//2 inputs
        syndrom[ 8] = in[ 4]^in[10];//2 inputs
        syndrom[ 9] = in[ 4]^in[11];//2 inputs
        syndrom[10] = in[ 5]^in[10];//2 inputs
        syndrom[11] = in[ 5]^in[11];//2 inputs
        syndrom[12] = in[ 6]^in[ 8];//2 inputs
        syndrom[13] = in[ 6]^in[ 9];//2 inputs
        syndrom[14] = in[ 7]^in[ 8];//2 inputs
        syndrom[15] = in[ 7]^in[ 9];//2 inputs
        hamming_code_32_16_f = syndrom;
    end
endfunction
wire [16-1:0] stored_data_edc = hamming_code_32_16_f(i_stored_data);
wire [16-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_16_min_delay (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [16-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [16-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_32_16_f
//Compute 16 bits Error Detection Code from a 16 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 4294967296 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[ 0]: x        x  x    (3 inputs)
//  syndrom[ 1]: x         xx     (3 inputs)
//  syndrom[ 2]: x         xx     (3 inputs)
//  syndrom[ 3]:  x      x    x   (3 inputs)
//  syndrom[ 4]:  x       xx      (3 inputs)
//  syndrom[ 5]:  x       x x     (3 inputs)
//  syndrom[ 6]:   x    x      x  (3 inputs)
//  syndrom[ 7]:   x     x   x    (3 inputs)
//  syndrom[ 8]:   x     x   x    (3 inputs)
//  syndrom[ 9]:    x  x        x (3 inputs)
//  syndrom[10]:    x   x     x   (3 inputs)
//  syndrom[11]:    x   x     x   (3 inputs)
//  syndrom[12]:     xx         x (3 inputs)
//  syndrom[13]:     xx         x (3 inputs)
//  syndrom[14]:     x x       x  (3 inputs)
//  syndrom[15]:      xx       x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 12 13 15)
//  input bit  6 used  3 times (syndrom bits 9 14 15)
//  input bit  7 used  3 times (syndrom bits 6 10 11)
//  input bit  8 used  3 times (syndrom bits 3 7 8)
//  input bit  9 used  3 times (syndrom bits 0 4 5)
//  input bit 10 used  3 times (syndrom bits 1 2 4)
//  input bit 11 used  3 times (syndrom bits 1 2 5)
//  input bit 12 used  3 times (syndrom bits 0 7 8)
//  input bit 13 used  3 times (syndrom bits 3 10 11)
//  input bit 14 used  3 times (syndrom bits 6 14 15)
//  input bit 15 used  3 times (syndrom bits 9 12 13)
function [16-1:0] extended_hamming_code_32_16_f;
    input [16-1:0] in;
    reg [16-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 9]^in[12];//3 inputs
        syndrom[ 1] = in[ 0]^in[10]^in[11];//3 inputs
        syndrom[ 2] = in[ 0]^in[10]^in[11];//3 inputs
        syndrom[ 3] = in[ 1]^in[ 8]^in[13];//3 inputs
        syndrom[ 4] = in[ 1]^in[ 9]^in[10];//3 inputs
        syndrom[ 5] = in[ 1]^in[ 9]^in[11];//3 inputs
        syndrom[ 6] = in[ 2]^in[ 7]^in[14];//3 inputs
        syndrom[ 7] = in[ 2]^in[ 8]^in[12];//3 inputs
        syndrom[ 8] = in[ 2]^in[ 8]^in[12];//3 inputs
        syndrom[ 9] = in[ 3]^in[ 6]^in[15];//3 inputs
        syndrom[10] = in[ 3]^in[ 7]^in[13];//3 inputs
        syndrom[11] = in[ 3]^in[ 7]^in[13];//3 inputs
        syndrom[12] = in[ 4]^in[ 5]^in[15];//3 inputs
        syndrom[13] = in[ 4]^in[ 5]^in[15];//3 inputs
        syndrom[14] = in[ 4]^in[ 6]^in[14];//3 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[14];//3 inputs
        extended_hamming_code_32_16_f = syndrom;
    end
endfunction
wire [16-1:0] stored_data_edc = extended_hamming_code_32_16_f(i_stored_data);
wire [16-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_16_min_delay (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [16-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [16-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [16-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_32_16_f
//Compute 16 bits Error Detection Code from a 16 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 4294967296 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[ 0]: x        x  x    (3 inputs)
//  syndrom[ 1]: x         xx     (3 inputs)
//  syndrom[ 2]: x         xx     (3 inputs)
//  syndrom[ 3]:  x      x    x   (3 inputs)
//  syndrom[ 4]:  x       xx      (3 inputs)
//  syndrom[ 5]:  x       x x     (3 inputs)
//  syndrom[ 6]:   x    x      x  (3 inputs)
//  syndrom[ 7]:   x     x   x    (3 inputs)
//  syndrom[ 8]:   x     x   x    (3 inputs)
//  syndrom[ 9]:    x  x        x (3 inputs)
//  syndrom[10]:    x   x     x   (3 inputs)
//  syndrom[11]:    x   x     x   (3 inputs)
//  syndrom[12]:     xx         x (3 inputs)
//  syndrom[13]:     xx         x (3 inputs)
//  syndrom[14]:     x x       x  (3 inputs)
//  syndrom[15]:      xx       x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 12 13 15)
//  input bit  6 used  3 times (syndrom bits 9 14 15)
//  input bit  7 used  3 times (syndrom bits 6 10 11)
//  input bit  8 used  3 times (syndrom bits 3 7 8)
//  input bit  9 used  3 times (syndrom bits 0 4 5)
//  input bit 10 used  3 times (syndrom bits 1 2 4)
//  input bit 11 used  3 times (syndrom bits 1 2 5)
//  input bit 12 used  3 times (syndrom bits 0 7 8)
//  input bit 13 used  3 times (syndrom bits 3 10 11)
//  input bit 14 used  3 times (syndrom bits 6 14 15)
//  input bit 15 used  3 times (syndrom bits 9 12 13)
function [16-1:0] extended_hamming_code_32_16_f;
    input [16-1:0] in;
    reg [16-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 9]^in[12];//3 inputs
        syndrom[ 1] = in[ 0]^in[10]^in[11];//3 inputs
        syndrom[ 2] = in[ 0]^in[10]^in[11];//3 inputs
        syndrom[ 3] = in[ 1]^in[ 8]^in[13];//3 inputs
        syndrom[ 4] = in[ 1]^in[ 9]^in[10];//3 inputs
        syndrom[ 5] = in[ 1]^in[ 9]^in[11];//3 inputs
        syndrom[ 6] = in[ 2]^in[ 7]^in[14];//3 inputs
        syndrom[ 7] = in[ 2]^in[ 8]^in[12];//3 inputs
        syndrom[ 8] = in[ 2]^in[ 8]^in[12];//3 inputs
        syndrom[ 9] = in[ 3]^in[ 6]^in[15];//3 inputs
        syndrom[10] = in[ 3]^in[ 7]^in[13];//3 inputs
        syndrom[11] = in[ 3]^in[ 7]^in[13];//3 inputs
        syndrom[12] = in[ 4]^in[ 5]^in[15];//3 inputs
        syndrom[13] = in[ 4]^in[ 5]^in[15];//3 inputs
        syndrom[14] = in[ 4]^in[ 6]^in[14];//3 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[14];//3 inputs
        extended_hamming_code_32_16_f = syndrom;
    end
endfunction
function [2+16-1:0] extended_hamming_code_32_16_f_correction_pattern_f;
    input [16-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [16-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {16{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			16'b0000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {16{1'b0}};
			end	
			16'b0000000000000111: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 0]=1'b1;
			end
			16'b0000000000111000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 1]=1'b1;
			end
			16'b0000000111000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 2]=1'b1;
			end
			16'b0000111000000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 3]=1'b1;
			end
			16'b0111000000000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 4]=1'b1;
			end
			16'b1011000000000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 5]=1'b1;
			end
			16'b1100001000000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 6]=1'b1;
			end
			16'b0000110001000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 7]=1'b1;
			end
			16'b0000000110001000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 8]=1'b1;
			end
			16'b0000000000110001: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 9]=1'b1;
			end
			16'b0000000000010110: begin
				correction_pattern = {16{1'b0}};correction_pattern[10]=1'b1;
			end
			16'b0000000000100110: begin
				correction_pattern = {16{1'b0}};correction_pattern[11]=1'b1;
			end
			16'b0000000110000001: begin
				correction_pattern = {16{1'b0}};correction_pattern[12]=1'b1;
			end
			16'b0000110000001000: begin
				correction_pattern = {16{1'b0}};correction_pattern[13]=1'b1;
			end
			16'b1100000001000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[14]=1'b1;
			end
			16'b0011001000000000: begin
				correction_pattern = {16{1'b0}};correction_pattern[15]=1'b1;
			end
			16'b0000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b1000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_32_16_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [16-1:0] stored_data_edc = extended_hamming_code_32_16_f(i_stored_data);
wire [16-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [16-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_32_16_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_20_min_delay (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [20-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [20-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_40_20_f
//Compute 20 bits Error Detection Code from a 20 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 1099511627776 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[ 0]: x                 x  (2 inputs)
//  syndrom[ 1]: x                  x (2 inputs)
//  syndrom[ 2]:  x                x  (2 inputs)
//  syndrom[ 3]:  x                 x (2 inputs)
//  syndrom[ 4]:   x             x    (2 inputs)
//  syndrom[ 5]:   x              x   (2 inputs)
//  syndrom[ 6]:    x            x    (2 inputs)
//  syndrom[ 7]:    x             x   (2 inputs)
//  syndrom[ 8]:     x         x      (2 inputs)
//  syndrom[ 9]:     x          x     (2 inputs)
//  syndrom[10]:      x        x      (2 inputs)
//  syndrom[11]:      x         x     (2 inputs)
//  syndrom[12]:       x     x        (2 inputs)
//  syndrom[13]:       x      x       (2 inputs)
//  syndrom[14]:        x    x        (2 inputs)
//  syndrom[15]:        x     x       (2 inputs)
//  syndrom[16]:         x x          (2 inputs)
//  syndrom[17]:         x  x         (2 inputs)
//  syndrom[18]:          xx          (2 inputs)
//  syndrom[19]:          x x         (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 16 18)
//  input bit 11 used  2 times (syndrom bits 17 19)
//  input bit 12 used  2 times (syndrom bits 12 14)
//  input bit 13 used  2 times (syndrom bits 13 15)
//  input bit 14 used  2 times (syndrom bits 8 10)
//  input bit 15 used  2 times (syndrom bits 9 11)
//  input bit 16 used  2 times (syndrom bits 4 6)
//  input bit 17 used  2 times (syndrom bits 5 7)
//  input bit 18 used  2 times (syndrom bits 0 2)
//  input bit 19 used  2 times (syndrom bits 1 3)
function [20-1:0] hamming_code_40_20_f;
    input [20-1:0] in;
    reg [20-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[18];//2 inputs
        syndrom[ 1] = in[ 0]^in[19];//2 inputs
        syndrom[ 2] = in[ 1]^in[18];//2 inputs
        syndrom[ 3] = in[ 1]^in[19];//2 inputs
        syndrom[ 4] = in[ 2]^in[16];//2 inputs
        syndrom[ 5] = in[ 2]^in[17];//2 inputs
        syndrom[ 6] = in[ 3]^in[16];//2 inputs
        syndrom[ 7] = in[ 3]^in[17];//2 inputs
        syndrom[ 8] = in[ 4]^in[14];//2 inputs
        syndrom[ 9] = in[ 4]^in[15];//2 inputs
        syndrom[10] = in[ 5]^in[14];//2 inputs
        syndrom[11] = in[ 5]^in[15];//2 inputs
        syndrom[12] = in[ 6]^in[12];//2 inputs
        syndrom[13] = in[ 6]^in[13];//2 inputs
        syndrom[14] = in[ 7]^in[12];//2 inputs
        syndrom[15] = in[ 7]^in[13];//2 inputs
        syndrom[16] = in[ 8]^in[10];//2 inputs
        syndrom[17] = in[ 8]^in[11];//2 inputs
        syndrom[18] = in[ 9]^in[10];//2 inputs
        syndrom[19] = in[ 9]^in[11];//2 inputs
        hamming_code_40_20_f = syndrom;
    end
endfunction
wire [20-1:0] stored_data_edc = hamming_code_40_20_f(i_stored_data);
wire [20-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_20_min_delay (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [20-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [20-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_40_20_f
//Compute 20 bits Error Detection Code from a 20 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 1099511627776 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[ 0]: x           xx       (3 inputs)
//  syndrom[ 1]: x           x x      (3 inputs)
//  syndrom[ 2]: x            xx      (3 inputs)
//  syndrom[ 3]:  x         x   x     (3 inputs)
//  syndrom[ 4]:  x         x   x     (3 inputs)
//  syndrom[ 5]:  x          xx       (3 inputs)
//  syndrom[ 6]:   x       x     x    (3 inputs)
//  syndrom[ 7]:   x       x     x    (3 inputs)
//  syndrom[ 8]:   x        x  x      (3 inputs)
//  syndrom[ 9]:    x     x       x   (3 inputs)
//  syndrom[10]:    x     x       x   (3 inputs)
//  syndrom[11]:    x      x    x     (3 inputs)
//  syndrom[12]:     x   x         x  (3 inputs)
//  syndrom[13]:     x   x         x  (3 inputs)
//  syndrom[14]:     x    x      x    (3 inputs)
//  syndrom[15]:      xx            x (3 inputs)
//  syndrom[16]:      x x           x (3 inputs)
//  syndrom[17]:      x  x        x   (3 inputs)
//  syndrom[18]:       xx          x  (3 inputs)
//  syndrom[19]:       xx           x (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 15 18 19)
//  input bit  7 used  3 times (syndrom bits 16 18 19)
//  input bit  8 used  3 times (syndrom bits 12 13 17)
//  input bit  9 used  3 times (syndrom bits 9 10 14)
//  input bit 10 used  3 times (syndrom bits 6 7 11)
//  input bit 11 used  3 times (syndrom bits 3 4 8)
//  input bit 12 used  3 times (syndrom bits 0 1 5)
//  input bit 13 used  3 times (syndrom bits 0 2 5)
//  input bit 14 used  3 times (syndrom bits 1 2 8)
//  input bit 15 used  3 times (syndrom bits 3 4 11)
//  input bit 16 used  3 times (syndrom bits 6 7 14)
//  input bit 17 used  3 times (syndrom bits 9 10 17)
//  input bit 18 used  3 times (syndrom bits 12 13 18)
//  input bit 19 used  3 times (syndrom bits 15 16 19)
function [20-1:0] extended_hamming_code_40_20_f;
    input [20-1:0] in;
    reg [20-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[12]^in[13];//3 inputs
        syndrom[ 1] = in[ 0]^in[12]^in[14];//3 inputs
        syndrom[ 2] = in[ 0]^in[13]^in[14];//3 inputs
        syndrom[ 3] = in[ 1]^in[11]^in[15];//3 inputs
        syndrom[ 4] = in[ 1]^in[11]^in[15];//3 inputs
        syndrom[ 5] = in[ 1]^in[12]^in[13];//3 inputs
        syndrom[ 6] = in[ 2]^in[10]^in[16];//3 inputs
        syndrom[ 7] = in[ 2]^in[10]^in[16];//3 inputs
        syndrom[ 8] = in[ 2]^in[11]^in[14];//3 inputs
        syndrom[ 9] = in[ 3]^in[ 9]^in[17];//3 inputs
        syndrom[10] = in[ 3]^in[ 9]^in[17];//3 inputs
        syndrom[11] = in[ 3]^in[10]^in[15];//3 inputs
        syndrom[12] = in[ 4]^in[ 8]^in[18];//3 inputs
        syndrom[13] = in[ 4]^in[ 8]^in[18];//3 inputs
        syndrom[14] = in[ 4]^in[ 9]^in[16];//3 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[19];//3 inputs
        syndrom[16] = in[ 5]^in[ 7]^in[19];//3 inputs
        syndrom[17] = in[ 5]^in[ 8]^in[17];//3 inputs
        syndrom[18] = in[ 6]^in[ 7]^in[18];//3 inputs
        syndrom[19] = in[ 6]^in[ 7]^in[19];//3 inputs
        extended_hamming_code_40_20_f = syndrom;
    end
endfunction
wire [20-1:0] stored_data_edc = extended_hamming_code_40_20_f(i_stored_data);
wire [20-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_20_min_delay (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [20-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [20-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [20-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_40_20_f
//Compute 20 bits Error Detection Code from a 20 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 1099511627776 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[ 0]: x           xx       (3 inputs)
//  syndrom[ 1]: x           x x      (3 inputs)
//  syndrom[ 2]: x            xx      (3 inputs)
//  syndrom[ 3]:  x         x   x     (3 inputs)
//  syndrom[ 4]:  x         x   x     (3 inputs)
//  syndrom[ 5]:  x          xx       (3 inputs)
//  syndrom[ 6]:   x       x     x    (3 inputs)
//  syndrom[ 7]:   x       x     x    (3 inputs)
//  syndrom[ 8]:   x        x  x      (3 inputs)
//  syndrom[ 9]:    x     x       x   (3 inputs)
//  syndrom[10]:    x     x       x   (3 inputs)
//  syndrom[11]:    x      x    x     (3 inputs)
//  syndrom[12]:     x   x         x  (3 inputs)
//  syndrom[13]:     x   x         x  (3 inputs)
//  syndrom[14]:     x    x      x    (3 inputs)
//  syndrom[15]:      xx            x (3 inputs)
//  syndrom[16]:      x x           x (3 inputs)
//  syndrom[17]:      x  x        x   (3 inputs)
//  syndrom[18]:       xx          x  (3 inputs)
//  syndrom[19]:       xx           x (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 15 18 19)
//  input bit  7 used  3 times (syndrom bits 16 18 19)
//  input bit  8 used  3 times (syndrom bits 12 13 17)
//  input bit  9 used  3 times (syndrom bits 9 10 14)
//  input bit 10 used  3 times (syndrom bits 6 7 11)
//  input bit 11 used  3 times (syndrom bits 3 4 8)
//  input bit 12 used  3 times (syndrom bits 0 1 5)
//  input bit 13 used  3 times (syndrom bits 0 2 5)
//  input bit 14 used  3 times (syndrom bits 1 2 8)
//  input bit 15 used  3 times (syndrom bits 3 4 11)
//  input bit 16 used  3 times (syndrom bits 6 7 14)
//  input bit 17 used  3 times (syndrom bits 9 10 17)
//  input bit 18 used  3 times (syndrom bits 12 13 18)
//  input bit 19 used  3 times (syndrom bits 15 16 19)
function [20-1:0] extended_hamming_code_40_20_f;
    input [20-1:0] in;
    reg [20-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[12]^in[13];//3 inputs
        syndrom[ 1] = in[ 0]^in[12]^in[14];//3 inputs
        syndrom[ 2] = in[ 0]^in[13]^in[14];//3 inputs
        syndrom[ 3] = in[ 1]^in[11]^in[15];//3 inputs
        syndrom[ 4] = in[ 1]^in[11]^in[15];//3 inputs
        syndrom[ 5] = in[ 1]^in[12]^in[13];//3 inputs
        syndrom[ 6] = in[ 2]^in[10]^in[16];//3 inputs
        syndrom[ 7] = in[ 2]^in[10]^in[16];//3 inputs
        syndrom[ 8] = in[ 2]^in[11]^in[14];//3 inputs
        syndrom[ 9] = in[ 3]^in[ 9]^in[17];//3 inputs
        syndrom[10] = in[ 3]^in[ 9]^in[17];//3 inputs
        syndrom[11] = in[ 3]^in[10]^in[15];//3 inputs
        syndrom[12] = in[ 4]^in[ 8]^in[18];//3 inputs
        syndrom[13] = in[ 4]^in[ 8]^in[18];//3 inputs
        syndrom[14] = in[ 4]^in[ 9]^in[16];//3 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[19];//3 inputs
        syndrom[16] = in[ 5]^in[ 7]^in[19];//3 inputs
        syndrom[17] = in[ 5]^in[ 8]^in[17];//3 inputs
        syndrom[18] = in[ 6]^in[ 7]^in[18];//3 inputs
        syndrom[19] = in[ 6]^in[ 7]^in[19];//3 inputs
        extended_hamming_code_40_20_f = syndrom;
    end
endfunction
function [2+20-1:0] extended_hamming_code_40_20_f_correction_pattern_f;
    input [20-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [20-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {20{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			20'b00000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {20{1'b0}};
			end	
			20'b00000000000000000111: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 0]=1'b1;
			end
			20'b00000000000000111000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 1]=1'b1;
			end
			20'b00000000000111000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 2]=1'b1;
			end
			20'b00000000111000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 3]=1'b1;
			end
			20'b00000111000000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 4]=1'b1;
			end
			20'b00111000000000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 5]=1'b1;
			end
			20'b11001000000000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 6]=1'b1;
			end
			20'b11010000000000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 7]=1'b1;
			end
			20'b00100011000000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 8]=1'b1;
			end
			20'b00000100011000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 9]=1'b1;
			end
			20'b00000000100011000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[10]=1'b1;
			end
			20'b00000000000100011000: begin
				correction_pattern = {20{1'b0}};correction_pattern[11]=1'b1;
			end
			20'b00000000000000100011: begin
				correction_pattern = {20{1'b0}};correction_pattern[12]=1'b1;
			end
			20'b00000000000000100101: begin
				correction_pattern = {20{1'b0}};correction_pattern[13]=1'b1;
			end
			20'b00000000000100000110: begin
				correction_pattern = {20{1'b0}};correction_pattern[14]=1'b1;
			end
			20'b00000000100000011000: begin
				correction_pattern = {20{1'b0}};correction_pattern[15]=1'b1;
			end
			20'b00000100000011000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[16]=1'b1;
			end
			20'b00100000011000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[17]=1'b1;
			end
			20'b01000011000000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[18]=1'b1;
			end
			20'b10011000000000000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[19]=1'b1;
			end
			20'b00000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b01000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b10000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_40_20_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [20-1:0] stored_data_edc = extended_hamming_code_40_20_f(i_stored_data);
wire [20-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [20-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_40_20_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_24_min_delay (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [24-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [24-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_48_24_f
//Compute 24 bits Error Detection Code from a 24 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 281474976710656 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[ 0]: x                     x  (2 inputs)
//  syndrom[ 1]: x                      x (2 inputs)
//  syndrom[ 2]:  x                    x  (2 inputs)
//  syndrom[ 3]:  x                     x (2 inputs)
//  syndrom[ 4]:   x                 x    (2 inputs)
//  syndrom[ 5]:   x                  x   (2 inputs)
//  syndrom[ 6]:    x                x    (2 inputs)
//  syndrom[ 7]:    x                 x   (2 inputs)
//  syndrom[ 8]:     x             x      (2 inputs)
//  syndrom[ 9]:     x              x     (2 inputs)
//  syndrom[10]:      x            x      (2 inputs)
//  syndrom[11]:      x             x     (2 inputs)
//  syndrom[12]:       x         x        (2 inputs)
//  syndrom[13]:       x          x       (2 inputs)
//  syndrom[14]:        x        x        (2 inputs)
//  syndrom[15]:        x         x       (2 inputs)
//  syndrom[16]:         x     x          (2 inputs)
//  syndrom[17]:         x      x         (2 inputs)
//  syndrom[18]:          x    x          (2 inputs)
//  syndrom[19]:          x     x         (2 inputs)
//  syndrom[20]:           x x            (2 inputs)
//  syndrom[21]:           x  x           (2 inputs)
//  syndrom[22]:            xx            (2 inputs)
//  syndrom[23]:            x x           (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 20 22)
//  input bit 13 used  2 times (syndrom bits 21 23)
//  input bit 14 used  2 times (syndrom bits 16 18)
//  input bit 15 used  2 times (syndrom bits 17 19)
//  input bit 16 used  2 times (syndrom bits 12 14)
//  input bit 17 used  2 times (syndrom bits 13 15)
//  input bit 18 used  2 times (syndrom bits 8 10)
//  input bit 19 used  2 times (syndrom bits 9 11)
//  input bit 20 used  2 times (syndrom bits 4 6)
//  input bit 21 used  2 times (syndrom bits 5 7)
//  input bit 22 used  2 times (syndrom bits 0 2)
//  input bit 23 used  2 times (syndrom bits 1 3)
function [24-1:0] hamming_code_48_24_f;
    input [24-1:0] in;
    reg [24-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[22];//2 inputs
        syndrom[ 1] = in[ 0]^in[23];//2 inputs
        syndrom[ 2] = in[ 1]^in[22];//2 inputs
        syndrom[ 3] = in[ 1]^in[23];//2 inputs
        syndrom[ 4] = in[ 2]^in[20];//2 inputs
        syndrom[ 5] = in[ 2]^in[21];//2 inputs
        syndrom[ 6] = in[ 3]^in[20];//2 inputs
        syndrom[ 7] = in[ 3]^in[21];//2 inputs
        syndrom[ 8] = in[ 4]^in[18];//2 inputs
        syndrom[ 9] = in[ 4]^in[19];//2 inputs
        syndrom[10] = in[ 5]^in[18];//2 inputs
        syndrom[11] = in[ 5]^in[19];//2 inputs
        syndrom[12] = in[ 6]^in[16];//2 inputs
        syndrom[13] = in[ 6]^in[17];//2 inputs
        syndrom[14] = in[ 7]^in[16];//2 inputs
        syndrom[15] = in[ 7]^in[17];//2 inputs
        syndrom[16] = in[ 8]^in[14];//2 inputs
        syndrom[17] = in[ 8]^in[15];//2 inputs
        syndrom[18] = in[ 9]^in[14];//2 inputs
        syndrom[19] = in[ 9]^in[15];//2 inputs
        syndrom[20] = in[10]^in[12];//2 inputs
        syndrom[21] = in[10]^in[13];//2 inputs
        syndrom[22] = in[11]^in[12];//2 inputs
        syndrom[23] = in[11]^in[13];//2 inputs
        hamming_code_48_24_f = syndrom;
    end
endfunction
wire [24-1:0] stored_data_edc = hamming_code_48_24_f(i_stored_data);
wire [24-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_24_min_delay (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [24-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [24-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_48_24_f
//Compute 24 bits Error Detection Code from a 24 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 281474976710656 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[ 0]: x             x  x       (3 inputs)
//  syndrom[ 1]: x              xx        (3 inputs)
//  syndrom[ 2]: x              x x       (3 inputs)
//  syndrom[ 3]:  x            x x        (3 inputs)
//  syndrom[ 4]:  x            x  x       (3 inputs)
//  syndrom[ 5]:  x             xx        (3 inputs)
//  syndrom[ 6]:   x         x      x     (3 inputs)
//  syndrom[ 7]:   x          x    x      (3 inputs)
//  syndrom[ 8]:   x          x     x     (3 inputs)
//  syndrom[ 9]:    x        x     x      (3 inputs)
//  syndrom[10]:    x        x      x     (3 inputs)
//  syndrom[11]:    x         x    x      (3 inputs)
//  syndrom[12]:     x     x          x   (3 inputs)
//  syndrom[13]:     x      x        x    (3 inputs)
//  syndrom[14]:     x      x         x   (3 inputs)
//  syndrom[15]:      x    x         x    (3 inputs)
//  syndrom[16]:      x    x          x   (3 inputs)
//  syndrom[17]:      x     x        x    (3 inputs)
//  syndrom[18]:       x x              x (3 inputs)
//  syndrom[19]:       x  x            x  (3 inputs)
//  syndrom[20]:       x  x             x (3 inputs)
//  syndrom[21]:        xx             x  (3 inputs)
//  syndrom[22]:        xx              x (3 inputs)
//  syndrom[23]:        x x            x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 18 21 22)
//  input bit  9 used  3 times (syndrom bits 19 20 23)
//  input bit 10 used  3 times (syndrom bits 12 15 16)
//  input bit 11 used  3 times (syndrom bits 13 14 17)
//  input bit 12 used  3 times (syndrom bits 6 9 10)
//  input bit 13 used  3 times (syndrom bits 7 8 11)
//  input bit 14 used  3 times (syndrom bits 0 3 4)
//  input bit 15 used  3 times (syndrom bits 1 2 5)
//  input bit 16 used  3 times (syndrom bits 1 3 5)
//  input bit 17 used  3 times (syndrom bits 0 2 4)
//  input bit 18 used  3 times (syndrom bits 7 9 11)
//  input bit 19 used  3 times (syndrom bits 6 8 10)
//  input bit 20 used  3 times (syndrom bits 13 15 17)
//  input bit 21 used  3 times (syndrom bits 12 14 16)
//  input bit 22 used  3 times (syndrom bits 19 21 23)
//  input bit 23 used  3 times (syndrom bits 18 20 22)
function [24-1:0] extended_hamming_code_48_24_f;
    input [24-1:0] in;
    reg [24-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[14]^in[17];//3 inputs
        syndrom[ 1] = in[ 0]^in[15]^in[16];//3 inputs
        syndrom[ 2] = in[ 0]^in[15]^in[17];//3 inputs
        syndrom[ 3] = in[ 1]^in[14]^in[16];//3 inputs
        syndrom[ 4] = in[ 1]^in[14]^in[17];//3 inputs
        syndrom[ 5] = in[ 1]^in[15]^in[16];//3 inputs
        syndrom[ 6] = in[ 2]^in[12]^in[19];//3 inputs
        syndrom[ 7] = in[ 2]^in[13]^in[18];//3 inputs
        syndrom[ 8] = in[ 2]^in[13]^in[19];//3 inputs
        syndrom[ 9] = in[ 3]^in[12]^in[18];//3 inputs
        syndrom[10] = in[ 3]^in[12]^in[19];//3 inputs
        syndrom[11] = in[ 3]^in[13]^in[18];//3 inputs
        syndrom[12] = in[ 4]^in[10]^in[21];//3 inputs
        syndrom[13] = in[ 4]^in[11]^in[20];//3 inputs
        syndrom[14] = in[ 4]^in[11]^in[21];//3 inputs
        syndrom[15] = in[ 5]^in[10]^in[20];//3 inputs
        syndrom[16] = in[ 5]^in[10]^in[21];//3 inputs
        syndrom[17] = in[ 5]^in[11]^in[20];//3 inputs
        syndrom[18] = in[ 6]^in[ 8]^in[23];//3 inputs
        syndrom[19] = in[ 6]^in[ 9]^in[22];//3 inputs
        syndrom[20] = in[ 6]^in[ 9]^in[23];//3 inputs
        syndrom[21] = in[ 7]^in[ 8]^in[22];//3 inputs
        syndrom[22] = in[ 7]^in[ 8]^in[23];//3 inputs
        syndrom[23] = in[ 7]^in[ 9]^in[22];//3 inputs
        extended_hamming_code_48_24_f = syndrom;
    end
endfunction
wire [24-1:0] stored_data_edc = extended_hamming_code_48_24_f(i_stored_data);
wire [24-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_24_min_delay (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [24-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [24-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [24-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_48_24_f
//Compute 24 bits Error Detection Code from a 24 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 281474976710656 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[ 0]: x             x  x       (3 inputs)
//  syndrom[ 1]: x              xx        (3 inputs)
//  syndrom[ 2]: x              x x       (3 inputs)
//  syndrom[ 3]:  x            x x        (3 inputs)
//  syndrom[ 4]:  x            x  x       (3 inputs)
//  syndrom[ 5]:  x             xx        (3 inputs)
//  syndrom[ 6]:   x         x      x     (3 inputs)
//  syndrom[ 7]:   x          x    x      (3 inputs)
//  syndrom[ 8]:   x          x     x     (3 inputs)
//  syndrom[ 9]:    x        x     x      (3 inputs)
//  syndrom[10]:    x        x      x     (3 inputs)
//  syndrom[11]:    x         x    x      (3 inputs)
//  syndrom[12]:     x     x          x   (3 inputs)
//  syndrom[13]:     x      x        x    (3 inputs)
//  syndrom[14]:     x      x         x   (3 inputs)
//  syndrom[15]:      x    x         x    (3 inputs)
//  syndrom[16]:      x    x          x   (3 inputs)
//  syndrom[17]:      x     x        x    (3 inputs)
//  syndrom[18]:       x x              x (3 inputs)
//  syndrom[19]:       x  x            x  (3 inputs)
//  syndrom[20]:       x  x             x (3 inputs)
//  syndrom[21]:        xx             x  (3 inputs)
//  syndrom[22]:        xx              x (3 inputs)
//  syndrom[23]:        x x            x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 18 21 22)
//  input bit  9 used  3 times (syndrom bits 19 20 23)
//  input bit 10 used  3 times (syndrom bits 12 15 16)
//  input bit 11 used  3 times (syndrom bits 13 14 17)
//  input bit 12 used  3 times (syndrom bits 6 9 10)
//  input bit 13 used  3 times (syndrom bits 7 8 11)
//  input bit 14 used  3 times (syndrom bits 0 3 4)
//  input bit 15 used  3 times (syndrom bits 1 2 5)
//  input bit 16 used  3 times (syndrom bits 1 3 5)
//  input bit 17 used  3 times (syndrom bits 0 2 4)
//  input bit 18 used  3 times (syndrom bits 7 9 11)
//  input bit 19 used  3 times (syndrom bits 6 8 10)
//  input bit 20 used  3 times (syndrom bits 13 15 17)
//  input bit 21 used  3 times (syndrom bits 12 14 16)
//  input bit 22 used  3 times (syndrom bits 19 21 23)
//  input bit 23 used  3 times (syndrom bits 18 20 22)
function [24-1:0] extended_hamming_code_48_24_f;
    input [24-1:0] in;
    reg [24-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[14]^in[17];//3 inputs
        syndrom[ 1] = in[ 0]^in[15]^in[16];//3 inputs
        syndrom[ 2] = in[ 0]^in[15]^in[17];//3 inputs
        syndrom[ 3] = in[ 1]^in[14]^in[16];//3 inputs
        syndrom[ 4] = in[ 1]^in[14]^in[17];//3 inputs
        syndrom[ 5] = in[ 1]^in[15]^in[16];//3 inputs
        syndrom[ 6] = in[ 2]^in[12]^in[19];//3 inputs
        syndrom[ 7] = in[ 2]^in[13]^in[18];//3 inputs
        syndrom[ 8] = in[ 2]^in[13]^in[19];//3 inputs
        syndrom[ 9] = in[ 3]^in[12]^in[18];//3 inputs
        syndrom[10] = in[ 3]^in[12]^in[19];//3 inputs
        syndrom[11] = in[ 3]^in[13]^in[18];//3 inputs
        syndrom[12] = in[ 4]^in[10]^in[21];//3 inputs
        syndrom[13] = in[ 4]^in[11]^in[20];//3 inputs
        syndrom[14] = in[ 4]^in[11]^in[21];//3 inputs
        syndrom[15] = in[ 5]^in[10]^in[20];//3 inputs
        syndrom[16] = in[ 5]^in[10]^in[21];//3 inputs
        syndrom[17] = in[ 5]^in[11]^in[20];//3 inputs
        syndrom[18] = in[ 6]^in[ 8]^in[23];//3 inputs
        syndrom[19] = in[ 6]^in[ 9]^in[22];//3 inputs
        syndrom[20] = in[ 6]^in[ 9]^in[23];//3 inputs
        syndrom[21] = in[ 7]^in[ 8]^in[22];//3 inputs
        syndrom[22] = in[ 7]^in[ 8]^in[23];//3 inputs
        syndrom[23] = in[ 7]^in[ 9]^in[22];//3 inputs
        extended_hamming_code_48_24_f = syndrom;
    end
endfunction
function [2+24-1:0] extended_hamming_code_48_24_f_correction_pattern_f;
    input [24-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [24-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {24{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			24'b000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {24{1'b0}};
			end	
			24'b000000000000000000000111: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 0]=1'b1;
			end
			24'b000000000000000000111000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 1]=1'b1;
			end
			24'b000000000000000111000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 2]=1'b1;
			end
			24'b000000000000111000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 3]=1'b1;
			end
			24'b000000000111000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 4]=1'b1;
			end
			24'b000000111000000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 5]=1'b1;
			end
			24'b000111000000000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 6]=1'b1;
			end
			24'b111000000000000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 7]=1'b1;
			end
			24'b011001000000000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 8]=1'b1;
			end
			24'b100110000000000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 9]=1'b1;
			end
			24'b000000011001000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[10]=1'b1;
			end
			24'b000000100110000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[11]=1'b1;
			end
			24'b000000000000011001000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[12]=1'b1;
			end
			24'b000000000000100110000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[13]=1'b1;
			end
			24'b000000000000000000011001: begin
				correction_pattern = {24{1'b0}};correction_pattern[14]=1'b1;
			end
			24'b000000000000000000100110: begin
				correction_pattern = {24{1'b0}};correction_pattern[15]=1'b1;
			end
			24'b000000000000000000101010: begin
				correction_pattern = {24{1'b0}};correction_pattern[16]=1'b1;
			end
			24'b000000000000000000010101: begin
				correction_pattern = {24{1'b0}};correction_pattern[17]=1'b1;
			end
			24'b000000000000101010000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[18]=1'b1;
			end
			24'b000000000000010101000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[19]=1'b1;
			end
			24'b000000101010000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[20]=1'b1;
			end
			24'b000000010101000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[21]=1'b1;
			end
			24'b101010000000000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[22]=1'b1;
			end
			24'b010101000000000000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[23]=1'b1;
			end
			24'b000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_48_24_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [24-1:0] stored_data_edc = extended_hamming_code_48_24_f(i_stored_data);
wire [24-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [24-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_48_24_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_32_min_delay (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [32-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [32-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_64_32_f
//Compute 32 bits Error Detection Code from a 32 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 18446744073709551616 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[ 0]: x                             x  (2 inputs)
//  syndrom[ 1]: x                              x (2 inputs)
//  syndrom[ 2]:  x                            x  (2 inputs)
//  syndrom[ 3]:  x                             x (2 inputs)
//  syndrom[ 4]:   x                         x    (2 inputs)
//  syndrom[ 5]:   x                          x   (2 inputs)
//  syndrom[ 6]:    x                        x    (2 inputs)
//  syndrom[ 7]:    x                         x   (2 inputs)
//  syndrom[ 8]:     x                     x      (2 inputs)
//  syndrom[ 9]:     x                      x     (2 inputs)
//  syndrom[10]:      x                    x      (2 inputs)
//  syndrom[11]:      x                     x     (2 inputs)
//  syndrom[12]:       x                 x        (2 inputs)
//  syndrom[13]:       x                  x       (2 inputs)
//  syndrom[14]:        x                x        (2 inputs)
//  syndrom[15]:        x                 x       (2 inputs)
//  syndrom[16]:         x             x          (2 inputs)
//  syndrom[17]:         x              x         (2 inputs)
//  syndrom[18]:          x            x          (2 inputs)
//  syndrom[19]:          x             x         (2 inputs)
//  syndrom[20]:           x         x            (2 inputs)
//  syndrom[21]:           x          x           (2 inputs)
//  syndrom[22]:            x        x            (2 inputs)
//  syndrom[23]:            x         x           (2 inputs)
//  syndrom[24]:             x     x              (2 inputs)
//  syndrom[25]:             x      x             (2 inputs)
//  syndrom[26]:              x    x              (2 inputs)
//  syndrom[27]:              x     x             (2 inputs)
//  syndrom[28]:               x x                (2 inputs)
//  syndrom[29]:               x  x               (2 inputs)
//  syndrom[30]:                xx                (2 inputs)
//  syndrom[31]:                x x               (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 28 30)
//  input bit 17 used  2 times (syndrom bits 29 31)
//  input bit 18 used  2 times (syndrom bits 24 26)
//  input bit 19 used  2 times (syndrom bits 25 27)
//  input bit 20 used  2 times (syndrom bits 20 22)
//  input bit 21 used  2 times (syndrom bits 21 23)
//  input bit 22 used  2 times (syndrom bits 16 18)
//  input bit 23 used  2 times (syndrom bits 17 19)
//  input bit 24 used  2 times (syndrom bits 12 14)
//  input bit 25 used  2 times (syndrom bits 13 15)
//  input bit 26 used  2 times (syndrom bits 8 10)
//  input bit 27 used  2 times (syndrom bits 9 11)
//  input bit 28 used  2 times (syndrom bits 4 6)
//  input bit 29 used  2 times (syndrom bits 5 7)
//  input bit 30 used  2 times (syndrom bits 0 2)
//  input bit 31 used  2 times (syndrom bits 1 3)
function [32-1:0] hamming_code_64_32_f;
    input [32-1:0] in;
    reg [32-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[30];//2 inputs
        syndrom[ 1] = in[ 0]^in[31];//2 inputs
        syndrom[ 2] = in[ 1]^in[30];//2 inputs
        syndrom[ 3] = in[ 1]^in[31];//2 inputs
        syndrom[ 4] = in[ 2]^in[28];//2 inputs
        syndrom[ 5] = in[ 2]^in[29];//2 inputs
        syndrom[ 6] = in[ 3]^in[28];//2 inputs
        syndrom[ 7] = in[ 3]^in[29];//2 inputs
        syndrom[ 8] = in[ 4]^in[26];//2 inputs
        syndrom[ 9] = in[ 4]^in[27];//2 inputs
        syndrom[10] = in[ 5]^in[26];//2 inputs
        syndrom[11] = in[ 5]^in[27];//2 inputs
        syndrom[12] = in[ 6]^in[24];//2 inputs
        syndrom[13] = in[ 6]^in[25];//2 inputs
        syndrom[14] = in[ 7]^in[24];//2 inputs
        syndrom[15] = in[ 7]^in[25];//2 inputs
        syndrom[16] = in[ 8]^in[22];//2 inputs
        syndrom[17] = in[ 8]^in[23];//2 inputs
        syndrom[18] = in[ 9]^in[22];//2 inputs
        syndrom[19] = in[ 9]^in[23];//2 inputs
        syndrom[20] = in[10]^in[20];//2 inputs
        syndrom[21] = in[10]^in[21];//2 inputs
        syndrom[22] = in[11]^in[20];//2 inputs
        syndrom[23] = in[11]^in[21];//2 inputs
        syndrom[24] = in[12]^in[18];//2 inputs
        syndrom[25] = in[12]^in[19];//2 inputs
        syndrom[26] = in[13]^in[18];//2 inputs
        syndrom[27] = in[13]^in[19];//2 inputs
        syndrom[28] = in[14]^in[16];//2 inputs
        syndrom[29] = in[14]^in[17];//2 inputs
        syndrom[30] = in[15]^in[16];//2 inputs
        syndrom[31] = in[15]^in[17];//2 inputs
        hamming_code_64_32_f = syndrom;
    end
endfunction
wire [32-1:0] stored_data_edc = hamming_code_64_32_f(i_stored_data);
wire [32-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_32_min_delay (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [32-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [32-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_64_32_f
//Compute 32 bits Error Detection Code from a 32 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 18446744073709551616 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[ 0]: x                   xx           (3 inputs)
//  syndrom[ 1]: x                   x x          (3 inputs)
//  syndrom[ 2]: x                    xx          (3 inputs)
//  syndrom[ 3]:  x                 x   x         (3 inputs)
//  syndrom[ 4]:  x                 x   x         (3 inputs)
//  syndrom[ 5]:  x                  xx           (3 inputs)
//  syndrom[ 6]:   x               x     x        (3 inputs)
//  syndrom[ 7]:   x               x     x        (3 inputs)
//  syndrom[ 8]:   x                x  x          (3 inputs)
//  syndrom[ 9]:    x             x       x       (3 inputs)
//  syndrom[10]:    x             x       x       (3 inputs)
//  syndrom[11]:    x              x    x         (3 inputs)
//  syndrom[12]:     x           x         x      (3 inputs)
//  syndrom[13]:     x           x         x      (3 inputs)
//  syndrom[14]:     x            x      x        (3 inputs)
//  syndrom[15]:      x         x           x     (3 inputs)
//  syndrom[16]:      x         x           x     (3 inputs)
//  syndrom[17]:      x          x        x       (3 inputs)
//  syndrom[18]:       x       x             x    (3 inputs)
//  syndrom[19]:       x       x             x    (3 inputs)
//  syndrom[20]:       x        x          x      (3 inputs)
//  syndrom[21]:        x     x               x   (3 inputs)
//  syndrom[22]:        x     x               x   (3 inputs)
//  syndrom[23]:        x      x            x     (3 inputs)
//  syndrom[24]:         x   x                 x  (3 inputs)
//  syndrom[25]:         x   x                 x  (3 inputs)
//  syndrom[26]:         x    x              x    (3 inputs)
//  syndrom[27]:          xx                    x (3 inputs)
//  syndrom[28]:          x x                   x (3 inputs)
//  syndrom[29]:          x  x                x   (3 inputs)
//  syndrom[30]:           xx                  x  (3 inputs)
//  syndrom[31]:           xx                   x (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 27 30 31)
//  input bit 11 used  3 times (syndrom bits 28 30 31)
//  input bit 12 used  3 times (syndrom bits 24 25 29)
//  input bit 13 used  3 times (syndrom bits 21 22 26)
//  input bit 14 used  3 times (syndrom bits 18 19 23)
//  input bit 15 used  3 times (syndrom bits 15 16 20)
//  input bit 16 used  3 times (syndrom bits 12 13 17)
//  input bit 17 used  3 times (syndrom bits 9 10 14)
//  input bit 18 used  3 times (syndrom bits 6 7 11)
//  input bit 19 used  3 times (syndrom bits 3 4 8)
//  input bit 20 used  3 times (syndrom bits 0 1 5)
//  input bit 21 used  3 times (syndrom bits 0 2 5)
//  input bit 22 used  3 times (syndrom bits 1 2 8)
//  input bit 23 used  3 times (syndrom bits 3 4 11)
//  input bit 24 used  3 times (syndrom bits 6 7 14)
//  input bit 25 used  3 times (syndrom bits 9 10 17)
//  input bit 26 used  3 times (syndrom bits 12 13 20)
//  input bit 27 used  3 times (syndrom bits 15 16 23)
//  input bit 28 used  3 times (syndrom bits 18 19 26)
//  input bit 29 used  3 times (syndrom bits 21 22 29)
//  input bit 30 used  3 times (syndrom bits 24 25 30)
//  input bit 31 used  3 times (syndrom bits 27 28 31)
function [32-1:0] extended_hamming_code_64_32_f;
    input [32-1:0] in;
    reg [32-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[20]^in[21];//3 inputs
        syndrom[ 1] = in[ 0]^in[20]^in[22];//3 inputs
        syndrom[ 2] = in[ 0]^in[21]^in[22];//3 inputs
        syndrom[ 3] = in[ 1]^in[19]^in[23];//3 inputs
        syndrom[ 4] = in[ 1]^in[19]^in[23];//3 inputs
        syndrom[ 5] = in[ 1]^in[20]^in[21];//3 inputs
        syndrom[ 6] = in[ 2]^in[18]^in[24];//3 inputs
        syndrom[ 7] = in[ 2]^in[18]^in[24];//3 inputs
        syndrom[ 8] = in[ 2]^in[19]^in[22];//3 inputs
        syndrom[ 9] = in[ 3]^in[17]^in[25];//3 inputs
        syndrom[10] = in[ 3]^in[17]^in[25];//3 inputs
        syndrom[11] = in[ 3]^in[18]^in[23];//3 inputs
        syndrom[12] = in[ 4]^in[16]^in[26];//3 inputs
        syndrom[13] = in[ 4]^in[16]^in[26];//3 inputs
        syndrom[14] = in[ 4]^in[17]^in[24];//3 inputs
        syndrom[15] = in[ 5]^in[15]^in[27];//3 inputs
        syndrom[16] = in[ 5]^in[15]^in[27];//3 inputs
        syndrom[17] = in[ 5]^in[16]^in[25];//3 inputs
        syndrom[18] = in[ 6]^in[14]^in[28];//3 inputs
        syndrom[19] = in[ 6]^in[14]^in[28];//3 inputs
        syndrom[20] = in[ 6]^in[15]^in[26];//3 inputs
        syndrom[21] = in[ 7]^in[13]^in[29];//3 inputs
        syndrom[22] = in[ 7]^in[13]^in[29];//3 inputs
        syndrom[23] = in[ 7]^in[14]^in[27];//3 inputs
        syndrom[24] = in[ 8]^in[12]^in[30];//3 inputs
        syndrom[25] = in[ 8]^in[12]^in[30];//3 inputs
        syndrom[26] = in[ 8]^in[13]^in[28];//3 inputs
        syndrom[27] = in[ 9]^in[10]^in[31];//3 inputs
        syndrom[28] = in[ 9]^in[11]^in[31];//3 inputs
        syndrom[29] = in[ 9]^in[12]^in[29];//3 inputs
        syndrom[30] = in[10]^in[11]^in[30];//3 inputs
        syndrom[31] = in[10]^in[11]^in[31];//3 inputs
        extended_hamming_code_64_32_f = syndrom;
    end
endfunction
wire [32-1:0] stored_data_edc = extended_hamming_code_64_32_f(i_stored_data);
wire [32-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_32_min_delay (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [32-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [32-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [32-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_64_32_f
//Compute 32 bits Error Detection Code from a 32 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 18446744073709551616 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[ 0]: x                   xx           (3 inputs)
//  syndrom[ 1]: x                   x x          (3 inputs)
//  syndrom[ 2]: x                    xx          (3 inputs)
//  syndrom[ 3]:  x                 x   x         (3 inputs)
//  syndrom[ 4]:  x                 x   x         (3 inputs)
//  syndrom[ 5]:  x                  xx           (3 inputs)
//  syndrom[ 6]:   x               x     x        (3 inputs)
//  syndrom[ 7]:   x               x     x        (3 inputs)
//  syndrom[ 8]:   x                x  x          (3 inputs)
//  syndrom[ 9]:    x             x       x       (3 inputs)
//  syndrom[10]:    x             x       x       (3 inputs)
//  syndrom[11]:    x              x    x         (3 inputs)
//  syndrom[12]:     x           x         x      (3 inputs)
//  syndrom[13]:     x           x         x      (3 inputs)
//  syndrom[14]:     x            x      x        (3 inputs)
//  syndrom[15]:      x         x           x     (3 inputs)
//  syndrom[16]:      x         x           x     (3 inputs)
//  syndrom[17]:      x          x        x       (3 inputs)
//  syndrom[18]:       x       x             x    (3 inputs)
//  syndrom[19]:       x       x             x    (3 inputs)
//  syndrom[20]:       x        x          x      (3 inputs)
//  syndrom[21]:        x     x               x   (3 inputs)
//  syndrom[22]:        x     x               x   (3 inputs)
//  syndrom[23]:        x      x            x     (3 inputs)
//  syndrom[24]:         x   x                 x  (3 inputs)
//  syndrom[25]:         x   x                 x  (3 inputs)
//  syndrom[26]:         x    x              x    (3 inputs)
//  syndrom[27]:          xx                    x (3 inputs)
//  syndrom[28]:          x x                   x (3 inputs)
//  syndrom[29]:          x  x                x   (3 inputs)
//  syndrom[30]:           xx                  x  (3 inputs)
//  syndrom[31]:           xx                   x (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 27 30 31)
//  input bit 11 used  3 times (syndrom bits 28 30 31)
//  input bit 12 used  3 times (syndrom bits 24 25 29)
//  input bit 13 used  3 times (syndrom bits 21 22 26)
//  input bit 14 used  3 times (syndrom bits 18 19 23)
//  input bit 15 used  3 times (syndrom bits 15 16 20)
//  input bit 16 used  3 times (syndrom bits 12 13 17)
//  input bit 17 used  3 times (syndrom bits 9 10 14)
//  input bit 18 used  3 times (syndrom bits 6 7 11)
//  input bit 19 used  3 times (syndrom bits 3 4 8)
//  input bit 20 used  3 times (syndrom bits 0 1 5)
//  input bit 21 used  3 times (syndrom bits 0 2 5)
//  input bit 22 used  3 times (syndrom bits 1 2 8)
//  input bit 23 used  3 times (syndrom bits 3 4 11)
//  input bit 24 used  3 times (syndrom bits 6 7 14)
//  input bit 25 used  3 times (syndrom bits 9 10 17)
//  input bit 26 used  3 times (syndrom bits 12 13 20)
//  input bit 27 used  3 times (syndrom bits 15 16 23)
//  input bit 28 used  3 times (syndrom bits 18 19 26)
//  input bit 29 used  3 times (syndrom bits 21 22 29)
//  input bit 30 used  3 times (syndrom bits 24 25 30)
//  input bit 31 used  3 times (syndrom bits 27 28 31)
function [32-1:0] extended_hamming_code_64_32_f;
    input [32-1:0] in;
    reg [32-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[20]^in[21];//3 inputs
        syndrom[ 1] = in[ 0]^in[20]^in[22];//3 inputs
        syndrom[ 2] = in[ 0]^in[21]^in[22];//3 inputs
        syndrom[ 3] = in[ 1]^in[19]^in[23];//3 inputs
        syndrom[ 4] = in[ 1]^in[19]^in[23];//3 inputs
        syndrom[ 5] = in[ 1]^in[20]^in[21];//3 inputs
        syndrom[ 6] = in[ 2]^in[18]^in[24];//3 inputs
        syndrom[ 7] = in[ 2]^in[18]^in[24];//3 inputs
        syndrom[ 8] = in[ 2]^in[19]^in[22];//3 inputs
        syndrom[ 9] = in[ 3]^in[17]^in[25];//3 inputs
        syndrom[10] = in[ 3]^in[17]^in[25];//3 inputs
        syndrom[11] = in[ 3]^in[18]^in[23];//3 inputs
        syndrom[12] = in[ 4]^in[16]^in[26];//3 inputs
        syndrom[13] = in[ 4]^in[16]^in[26];//3 inputs
        syndrom[14] = in[ 4]^in[17]^in[24];//3 inputs
        syndrom[15] = in[ 5]^in[15]^in[27];//3 inputs
        syndrom[16] = in[ 5]^in[15]^in[27];//3 inputs
        syndrom[17] = in[ 5]^in[16]^in[25];//3 inputs
        syndrom[18] = in[ 6]^in[14]^in[28];//3 inputs
        syndrom[19] = in[ 6]^in[14]^in[28];//3 inputs
        syndrom[20] = in[ 6]^in[15]^in[26];//3 inputs
        syndrom[21] = in[ 7]^in[13]^in[29];//3 inputs
        syndrom[22] = in[ 7]^in[13]^in[29];//3 inputs
        syndrom[23] = in[ 7]^in[14]^in[27];//3 inputs
        syndrom[24] = in[ 8]^in[12]^in[30];//3 inputs
        syndrom[25] = in[ 8]^in[12]^in[30];//3 inputs
        syndrom[26] = in[ 8]^in[13]^in[28];//3 inputs
        syndrom[27] = in[ 9]^in[10]^in[31];//3 inputs
        syndrom[28] = in[ 9]^in[11]^in[31];//3 inputs
        syndrom[29] = in[ 9]^in[12]^in[29];//3 inputs
        syndrom[30] = in[10]^in[11]^in[30];//3 inputs
        syndrom[31] = in[10]^in[11]^in[31];//3 inputs
        extended_hamming_code_64_32_f = syndrom;
    end
endfunction
function [2+32-1:0] extended_hamming_code_64_32_f_correction_pattern_f;
    input [32-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [32-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {32{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			32'b00000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {32{1'b0}};
			end	
			32'b00000000000000000000000000000111: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 0]=1'b1;
			end
			32'b00000000000000000000000000111000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 1]=1'b1;
			end
			32'b00000000000000000000000111000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 2]=1'b1;
			end
			32'b00000000000000000000111000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 3]=1'b1;
			end
			32'b00000000000000000111000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 4]=1'b1;
			end
			32'b00000000000000111000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 5]=1'b1;
			end
			32'b00000000000111000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 6]=1'b1;
			end
			32'b00000000111000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 7]=1'b1;
			end
			32'b00000111000000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 8]=1'b1;
			end
			32'b00111000000000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 9]=1'b1;
			end
			32'b11001000000000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[10]=1'b1;
			end
			32'b11010000000000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[11]=1'b1;
			end
			32'b00100011000000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[12]=1'b1;
			end
			32'b00000100011000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[13]=1'b1;
			end
			32'b00000000100011000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[14]=1'b1;
			end
			32'b00000000000100011000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[15]=1'b1;
			end
			32'b00000000000000100011000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[16]=1'b1;
			end
			32'b00000000000000000100011000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[17]=1'b1;
			end
			32'b00000000000000000000100011000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[18]=1'b1;
			end
			32'b00000000000000000000000100011000: begin
				correction_pattern = {32{1'b0}};correction_pattern[19]=1'b1;
			end
			32'b00000000000000000000000000100011: begin
				correction_pattern = {32{1'b0}};correction_pattern[20]=1'b1;
			end
			32'b00000000000000000000000000100101: begin
				correction_pattern = {32{1'b0}};correction_pattern[21]=1'b1;
			end
			32'b00000000000000000000000100000110: begin
				correction_pattern = {32{1'b0}};correction_pattern[22]=1'b1;
			end
			32'b00000000000000000000100000011000: begin
				correction_pattern = {32{1'b0}};correction_pattern[23]=1'b1;
			end
			32'b00000000000000000100000011000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[24]=1'b1;
			end
			32'b00000000000000100000011000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[25]=1'b1;
			end
			32'b00000000000100000011000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[26]=1'b1;
			end
			32'b00000000100000011000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[27]=1'b1;
			end
			32'b00000100000011000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[28]=1'b1;
			end
			32'b00100000011000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[29]=1'b1;
			end
			32'b01000011000000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[30]=1'b1;
			end
			32'b10011000000000000000000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[31]=1'b1;
			end
			32'b00000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b01000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b10000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_64_32_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [32-1:0] stored_data_edc = extended_hamming_code_64_32_f(i_stored_data);
wire [32-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [32-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_64_32_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_36_min_delay (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [36-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [36-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_72_36_f
//Compute 36 bits Error Detection Code from a 36 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[ 0]: x                                 x  (2 inputs)
//  syndrom[ 1]: x                                  x (2 inputs)
//  syndrom[ 2]:  x                                x  (2 inputs)
//  syndrom[ 3]:  x                                 x (2 inputs)
//  syndrom[ 4]:   x                             x    (2 inputs)
//  syndrom[ 5]:   x                              x   (2 inputs)
//  syndrom[ 6]:    x                            x    (2 inputs)
//  syndrom[ 7]:    x                             x   (2 inputs)
//  syndrom[ 8]:     x                         x      (2 inputs)
//  syndrom[ 9]:     x                          x     (2 inputs)
//  syndrom[10]:      x                        x      (2 inputs)
//  syndrom[11]:      x                         x     (2 inputs)
//  syndrom[12]:       x                     x        (2 inputs)
//  syndrom[13]:       x                      x       (2 inputs)
//  syndrom[14]:        x                    x        (2 inputs)
//  syndrom[15]:        x                     x       (2 inputs)
//  syndrom[16]:         x                 x          (2 inputs)
//  syndrom[17]:         x                  x         (2 inputs)
//  syndrom[18]:          x                x          (2 inputs)
//  syndrom[19]:          x                 x         (2 inputs)
//  syndrom[20]:           x             x            (2 inputs)
//  syndrom[21]:           x              x           (2 inputs)
//  syndrom[22]:            x            x            (2 inputs)
//  syndrom[23]:            x             x           (2 inputs)
//  syndrom[24]:             x         x              (2 inputs)
//  syndrom[25]:             x          x             (2 inputs)
//  syndrom[26]:              x        x              (2 inputs)
//  syndrom[27]:              x         x             (2 inputs)
//  syndrom[28]:               x     x                (2 inputs)
//  syndrom[29]:               x      x               (2 inputs)
//  syndrom[30]:                x    x                (2 inputs)
//  syndrom[31]:                x     x               (2 inputs)
//  syndrom[32]:                 x x                  (2 inputs)
//  syndrom[33]:                 x  x                 (2 inputs)
//  syndrom[34]:                  xx                  (2 inputs)
//  syndrom[35]:                  x x                 (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 32 33)
//  input bit 17 used  2 times (syndrom bits 34 35)
//  input bit 18 used  2 times (syndrom bits 32 34)
//  input bit 19 used  2 times (syndrom bits 33 35)
//  input bit 20 used  2 times (syndrom bits 28 30)
//  input bit 21 used  2 times (syndrom bits 29 31)
//  input bit 22 used  2 times (syndrom bits 24 26)
//  input bit 23 used  2 times (syndrom bits 25 27)
//  input bit 24 used  2 times (syndrom bits 20 22)
//  input bit 25 used  2 times (syndrom bits 21 23)
//  input bit 26 used  2 times (syndrom bits 16 18)
//  input bit 27 used  2 times (syndrom bits 17 19)
//  input bit 28 used  2 times (syndrom bits 12 14)
//  input bit 29 used  2 times (syndrom bits 13 15)
//  input bit 30 used  2 times (syndrom bits 8 10)
//  input bit 31 used  2 times (syndrom bits 9 11)
//  input bit 32 used  2 times (syndrom bits 4 6)
//  input bit 33 used  2 times (syndrom bits 5 7)
//  input bit 34 used  2 times (syndrom bits 0 2)
//  input bit 35 used  2 times (syndrom bits 1 3)
function [36-1:0] hamming_code_72_36_f;
    input [36-1:0] in;
    reg [36-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[34];//2 inputs
        syndrom[ 1] = in[ 0]^in[35];//2 inputs
        syndrom[ 2] = in[ 1]^in[34];//2 inputs
        syndrom[ 3] = in[ 1]^in[35];//2 inputs
        syndrom[ 4] = in[ 2]^in[32];//2 inputs
        syndrom[ 5] = in[ 2]^in[33];//2 inputs
        syndrom[ 6] = in[ 3]^in[32];//2 inputs
        syndrom[ 7] = in[ 3]^in[33];//2 inputs
        syndrom[ 8] = in[ 4]^in[30];//2 inputs
        syndrom[ 9] = in[ 4]^in[31];//2 inputs
        syndrom[10] = in[ 5]^in[30];//2 inputs
        syndrom[11] = in[ 5]^in[31];//2 inputs
        syndrom[12] = in[ 6]^in[28];//2 inputs
        syndrom[13] = in[ 6]^in[29];//2 inputs
        syndrom[14] = in[ 7]^in[28];//2 inputs
        syndrom[15] = in[ 7]^in[29];//2 inputs
        syndrom[16] = in[ 8]^in[26];//2 inputs
        syndrom[17] = in[ 8]^in[27];//2 inputs
        syndrom[18] = in[ 9]^in[26];//2 inputs
        syndrom[19] = in[ 9]^in[27];//2 inputs
        syndrom[20] = in[10]^in[24];//2 inputs
        syndrom[21] = in[10]^in[25];//2 inputs
        syndrom[22] = in[11]^in[24];//2 inputs
        syndrom[23] = in[11]^in[25];//2 inputs
        syndrom[24] = in[12]^in[22];//2 inputs
        syndrom[25] = in[12]^in[23];//2 inputs
        syndrom[26] = in[13]^in[22];//2 inputs
        syndrom[27] = in[13]^in[23];//2 inputs
        syndrom[28] = in[14]^in[20];//2 inputs
        syndrom[29] = in[14]^in[21];//2 inputs
        syndrom[30] = in[15]^in[20];//2 inputs
        syndrom[31] = in[15]^in[21];//2 inputs
        syndrom[32] = in[16]^in[18];//2 inputs
        syndrom[33] = in[16]^in[19];//2 inputs
        syndrom[34] = in[17]^in[18];//2 inputs
        syndrom[35] = in[17]^in[19];//2 inputs
        hamming_code_72_36_f = syndrom;
    end
endfunction
wire [36-1:0] stored_data_edc = hamming_code_72_36_f(i_stored_data);
wire [36-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_36_min_delay (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [36-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [36-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_72_36_f
//Compute 36 bits Error Detection Code from a 36 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[ 0]: x                     x  x           (3 inputs)
//  syndrom[ 1]: x                      xx            (3 inputs)
//  syndrom[ 2]: x                      x x           (3 inputs)
//  syndrom[ 3]:  x                    x x            (3 inputs)
//  syndrom[ 4]:  x                    x  x           (3 inputs)
//  syndrom[ 5]:  x                     xx            (3 inputs)
//  syndrom[ 6]:   x                 x      x         (3 inputs)
//  syndrom[ 7]:   x                  x    x          (3 inputs)
//  syndrom[ 8]:   x                  x     x         (3 inputs)
//  syndrom[ 9]:    x                x     x          (3 inputs)
//  syndrom[10]:    x                x      x         (3 inputs)
//  syndrom[11]:    x                 x    x          (3 inputs)
//  syndrom[12]:     x             x          x       (3 inputs)
//  syndrom[13]:     x              x        x        (3 inputs)
//  syndrom[14]:     x              x         x       (3 inputs)
//  syndrom[15]:      x            x         x        (3 inputs)
//  syndrom[16]:      x            x          x       (3 inputs)
//  syndrom[17]:      x             x        x        (3 inputs)
//  syndrom[18]:       x         x              x     (3 inputs)
//  syndrom[19]:       x          x            x      (3 inputs)
//  syndrom[20]:       x          x             x     (3 inputs)
//  syndrom[21]:        x        x             x      (3 inputs)
//  syndrom[22]:        x        x              x     (3 inputs)
//  syndrom[23]:        x         x            x      (3 inputs)
//  syndrom[24]:         x     x                  x   (3 inputs)
//  syndrom[25]:         x      x                x    (3 inputs)
//  syndrom[26]:         x      x                 x   (3 inputs)
//  syndrom[27]:          x    x                 x    (3 inputs)
//  syndrom[28]:          x    x                  x   (3 inputs)
//  syndrom[29]:          x     x                x    (3 inputs)
//  syndrom[30]:           x x                      x (3 inputs)
//  syndrom[31]:           x  x                    x  (3 inputs)
//  syndrom[32]:           x  x                     x (3 inputs)
//  syndrom[33]:            xx                     x  (3 inputs)
//  syndrom[34]:            xx                      x (3 inputs)
//  syndrom[35]:            x x                    x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 30 33 34)
//  input bit 13 used  3 times (syndrom bits 31 32 35)
//  input bit 14 used  3 times (syndrom bits 24 27 28)
//  input bit 15 used  3 times (syndrom bits 25 26 29)
//  input bit 16 used  3 times (syndrom bits 18 21 22)
//  input bit 17 used  3 times (syndrom bits 19 20 23)
//  input bit 18 used  3 times (syndrom bits 12 15 16)
//  input bit 19 used  3 times (syndrom bits 13 14 17)
//  input bit 20 used  3 times (syndrom bits 6 9 10)
//  input bit 21 used  3 times (syndrom bits 7 8 11)
//  input bit 22 used  3 times (syndrom bits 0 3 4)
//  input bit 23 used  3 times (syndrom bits 1 2 5)
//  input bit 24 used  3 times (syndrom bits 1 3 5)
//  input bit 25 used  3 times (syndrom bits 0 2 4)
//  input bit 26 used  3 times (syndrom bits 7 9 11)
//  input bit 27 used  3 times (syndrom bits 6 8 10)
//  input bit 28 used  3 times (syndrom bits 13 15 17)
//  input bit 29 used  3 times (syndrom bits 12 14 16)
//  input bit 30 used  3 times (syndrom bits 19 21 23)
//  input bit 31 used  3 times (syndrom bits 18 20 22)
//  input bit 32 used  3 times (syndrom bits 25 27 29)
//  input bit 33 used  3 times (syndrom bits 24 26 28)
//  input bit 34 used  3 times (syndrom bits 31 33 35)
//  input bit 35 used  3 times (syndrom bits 30 32 34)
function [36-1:0] extended_hamming_code_72_36_f;
    input [36-1:0] in;
    reg [36-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[22]^in[25];//3 inputs
        syndrom[ 1] = in[ 0]^in[23]^in[24];//3 inputs
        syndrom[ 2] = in[ 0]^in[23]^in[25];//3 inputs
        syndrom[ 3] = in[ 1]^in[22]^in[24];//3 inputs
        syndrom[ 4] = in[ 1]^in[22]^in[25];//3 inputs
        syndrom[ 5] = in[ 1]^in[23]^in[24];//3 inputs
        syndrom[ 6] = in[ 2]^in[20]^in[27];//3 inputs
        syndrom[ 7] = in[ 2]^in[21]^in[26];//3 inputs
        syndrom[ 8] = in[ 2]^in[21]^in[27];//3 inputs
        syndrom[ 9] = in[ 3]^in[20]^in[26];//3 inputs
        syndrom[10] = in[ 3]^in[20]^in[27];//3 inputs
        syndrom[11] = in[ 3]^in[21]^in[26];//3 inputs
        syndrom[12] = in[ 4]^in[18]^in[29];//3 inputs
        syndrom[13] = in[ 4]^in[19]^in[28];//3 inputs
        syndrom[14] = in[ 4]^in[19]^in[29];//3 inputs
        syndrom[15] = in[ 5]^in[18]^in[28];//3 inputs
        syndrom[16] = in[ 5]^in[18]^in[29];//3 inputs
        syndrom[17] = in[ 5]^in[19]^in[28];//3 inputs
        syndrom[18] = in[ 6]^in[16]^in[31];//3 inputs
        syndrom[19] = in[ 6]^in[17]^in[30];//3 inputs
        syndrom[20] = in[ 6]^in[17]^in[31];//3 inputs
        syndrom[21] = in[ 7]^in[16]^in[30];//3 inputs
        syndrom[22] = in[ 7]^in[16]^in[31];//3 inputs
        syndrom[23] = in[ 7]^in[17]^in[30];//3 inputs
        syndrom[24] = in[ 8]^in[14]^in[33];//3 inputs
        syndrom[25] = in[ 8]^in[15]^in[32];//3 inputs
        syndrom[26] = in[ 8]^in[15]^in[33];//3 inputs
        syndrom[27] = in[ 9]^in[14]^in[32];//3 inputs
        syndrom[28] = in[ 9]^in[14]^in[33];//3 inputs
        syndrom[29] = in[ 9]^in[15]^in[32];//3 inputs
        syndrom[30] = in[10]^in[12]^in[35];//3 inputs
        syndrom[31] = in[10]^in[13]^in[34];//3 inputs
        syndrom[32] = in[10]^in[13]^in[35];//3 inputs
        syndrom[33] = in[11]^in[12]^in[34];//3 inputs
        syndrom[34] = in[11]^in[12]^in[35];//3 inputs
        syndrom[35] = in[11]^in[13]^in[34];//3 inputs
        extended_hamming_code_72_36_f = syndrom;
    end
endfunction
wire [36-1:0] stored_data_edc = extended_hamming_code_72_36_f(i_stored_data);
wire [36-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_36_min_delay (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [36-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [36-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [36-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_72_36_f
//Compute 36 bits Error Detection Code from a 36 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[ 0]: x                     x  x           (3 inputs)
//  syndrom[ 1]: x                      xx            (3 inputs)
//  syndrom[ 2]: x                      x x           (3 inputs)
//  syndrom[ 3]:  x                    x x            (3 inputs)
//  syndrom[ 4]:  x                    x  x           (3 inputs)
//  syndrom[ 5]:  x                     xx            (3 inputs)
//  syndrom[ 6]:   x                 x      x         (3 inputs)
//  syndrom[ 7]:   x                  x    x          (3 inputs)
//  syndrom[ 8]:   x                  x     x         (3 inputs)
//  syndrom[ 9]:    x                x     x          (3 inputs)
//  syndrom[10]:    x                x      x         (3 inputs)
//  syndrom[11]:    x                 x    x          (3 inputs)
//  syndrom[12]:     x             x          x       (3 inputs)
//  syndrom[13]:     x              x        x        (3 inputs)
//  syndrom[14]:     x              x         x       (3 inputs)
//  syndrom[15]:      x            x         x        (3 inputs)
//  syndrom[16]:      x            x          x       (3 inputs)
//  syndrom[17]:      x             x        x        (3 inputs)
//  syndrom[18]:       x         x              x     (3 inputs)
//  syndrom[19]:       x          x            x      (3 inputs)
//  syndrom[20]:       x          x             x     (3 inputs)
//  syndrom[21]:        x        x             x      (3 inputs)
//  syndrom[22]:        x        x              x     (3 inputs)
//  syndrom[23]:        x         x            x      (3 inputs)
//  syndrom[24]:         x     x                  x   (3 inputs)
//  syndrom[25]:         x      x                x    (3 inputs)
//  syndrom[26]:         x      x                 x   (3 inputs)
//  syndrom[27]:          x    x                 x    (3 inputs)
//  syndrom[28]:          x    x                  x   (3 inputs)
//  syndrom[29]:          x     x                x    (3 inputs)
//  syndrom[30]:           x x                      x (3 inputs)
//  syndrom[31]:           x  x                    x  (3 inputs)
//  syndrom[32]:           x  x                     x (3 inputs)
//  syndrom[33]:            xx                     x  (3 inputs)
//  syndrom[34]:            xx                      x (3 inputs)
//  syndrom[35]:            x x                    x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 30 33 34)
//  input bit 13 used  3 times (syndrom bits 31 32 35)
//  input bit 14 used  3 times (syndrom bits 24 27 28)
//  input bit 15 used  3 times (syndrom bits 25 26 29)
//  input bit 16 used  3 times (syndrom bits 18 21 22)
//  input bit 17 used  3 times (syndrom bits 19 20 23)
//  input bit 18 used  3 times (syndrom bits 12 15 16)
//  input bit 19 used  3 times (syndrom bits 13 14 17)
//  input bit 20 used  3 times (syndrom bits 6 9 10)
//  input bit 21 used  3 times (syndrom bits 7 8 11)
//  input bit 22 used  3 times (syndrom bits 0 3 4)
//  input bit 23 used  3 times (syndrom bits 1 2 5)
//  input bit 24 used  3 times (syndrom bits 1 3 5)
//  input bit 25 used  3 times (syndrom bits 0 2 4)
//  input bit 26 used  3 times (syndrom bits 7 9 11)
//  input bit 27 used  3 times (syndrom bits 6 8 10)
//  input bit 28 used  3 times (syndrom bits 13 15 17)
//  input bit 29 used  3 times (syndrom bits 12 14 16)
//  input bit 30 used  3 times (syndrom bits 19 21 23)
//  input bit 31 used  3 times (syndrom bits 18 20 22)
//  input bit 32 used  3 times (syndrom bits 25 27 29)
//  input bit 33 used  3 times (syndrom bits 24 26 28)
//  input bit 34 used  3 times (syndrom bits 31 33 35)
//  input bit 35 used  3 times (syndrom bits 30 32 34)
function [36-1:0] extended_hamming_code_72_36_f;
    input [36-1:0] in;
    reg [36-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[22]^in[25];//3 inputs
        syndrom[ 1] = in[ 0]^in[23]^in[24];//3 inputs
        syndrom[ 2] = in[ 0]^in[23]^in[25];//3 inputs
        syndrom[ 3] = in[ 1]^in[22]^in[24];//3 inputs
        syndrom[ 4] = in[ 1]^in[22]^in[25];//3 inputs
        syndrom[ 5] = in[ 1]^in[23]^in[24];//3 inputs
        syndrom[ 6] = in[ 2]^in[20]^in[27];//3 inputs
        syndrom[ 7] = in[ 2]^in[21]^in[26];//3 inputs
        syndrom[ 8] = in[ 2]^in[21]^in[27];//3 inputs
        syndrom[ 9] = in[ 3]^in[20]^in[26];//3 inputs
        syndrom[10] = in[ 3]^in[20]^in[27];//3 inputs
        syndrom[11] = in[ 3]^in[21]^in[26];//3 inputs
        syndrom[12] = in[ 4]^in[18]^in[29];//3 inputs
        syndrom[13] = in[ 4]^in[19]^in[28];//3 inputs
        syndrom[14] = in[ 4]^in[19]^in[29];//3 inputs
        syndrom[15] = in[ 5]^in[18]^in[28];//3 inputs
        syndrom[16] = in[ 5]^in[18]^in[29];//3 inputs
        syndrom[17] = in[ 5]^in[19]^in[28];//3 inputs
        syndrom[18] = in[ 6]^in[16]^in[31];//3 inputs
        syndrom[19] = in[ 6]^in[17]^in[30];//3 inputs
        syndrom[20] = in[ 6]^in[17]^in[31];//3 inputs
        syndrom[21] = in[ 7]^in[16]^in[30];//3 inputs
        syndrom[22] = in[ 7]^in[16]^in[31];//3 inputs
        syndrom[23] = in[ 7]^in[17]^in[30];//3 inputs
        syndrom[24] = in[ 8]^in[14]^in[33];//3 inputs
        syndrom[25] = in[ 8]^in[15]^in[32];//3 inputs
        syndrom[26] = in[ 8]^in[15]^in[33];//3 inputs
        syndrom[27] = in[ 9]^in[14]^in[32];//3 inputs
        syndrom[28] = in[ 9]^in[14]^in[33];//3 inputs
        syndrom[29] = in[ 9]^in[15]^in[32];//3 inputs
        syndrom[30] = in[10]^in[12]^in[35];//3 inputs
        syndrom[31] = in[10]^in[13]^in[34];//3 inputs
        syndrom[32] = in[10]^in[13]^in[35];//3 inputs
        syndrom[33] = in[11]^in[12]^in[34];//3 inputs
        syndrom[34] = in[11]^in[12]^in[35];//3 inputs
        syndrom[35] = in[11]^in[13]^in[34];//3 inputs
        extended_hamming_code_72_36_f = syndrom;
    end
endfunction
function [2+36-1:0] extended_hamming_code_72_36_f_correction_pattern_f;
    input [36-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [36-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {36{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			36'b000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {36{1'b0}};
			end	
			36'b000000000000000000000000000000000111: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 0]=1'b1;
			end
			36'b000000000000000000000000000000111000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 1]=1'b1;
			end
			36'b000000000000000000000000000111000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 2]=1'b1;
			end
			36'b000000000000000000000000111000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 3]=1'b1;
			end
			36'b000000000000000000000111000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 4]=1'b1;
			end
			36'b000000000000000000111000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 5]=1'b1;
			end
			36'b000000000000000111000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 6]=1'b1;
			end
			36'b000000000000111000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 7]=1'b1;
			end
			36'b000000000111000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 8]=1'b1;
			end
			36'b000000111000000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 9]=1'b1;
			end
			36'b000111000000000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[10]=1'b1;
			end
			36'b111000000000000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[11]=1'b1;
			end
			36'b011001000000000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[12]=1'b1;
			end
			36'b100110000000000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[13]=1'b1;
			end
			36'b000000011001000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[14]=1'b1;
			end
			36'b000000100110000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[15]=1'b1;
			end
			36'b000000000000011001000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[16]=1'b1;
			end
			36'b000000000000100110000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[17]=1'b1;
			end
			36'b000000000000000000011001000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[18]=1'b1;
			end
			36'b000000000000000000100110000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[19]=1'b1;
			end
			36'b000000000000000000000000011001000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[20]=1'b1;
			end
			36'b000000000000000000000000100110000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[21]=1'b1;
			end
			36'b000000000000000000000000000000011001: begin
				correction_pattern = {36{1'b0}};correction_pattern[22]=1'b1;
			end
			36'b000000000000000000000000000000100110: begin
				correction_pattern = {36{1'b0}};correction_pattern[23]=1'b1;
			end
			36'b000000000000000000000000000000101010: begin
				correction_pattern = {36{1'b0}};correction_pattern[24]=1'b1;
			end
			36'b000000000000000000000000000000010101: begin
				correction_pattern = {36{1'b0}};correction_pattern[25]=1'b1;
			end
			36'b000000000000000000000000101010000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[26]=1'b1;
			end
			36'b000000000000000000000000010101000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[27]=1'b1;
			end
			36'b000000000000000000101010000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[28]=1'b1;
			end
			36'b000000000000000000010101000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[29]=1'b1;
			end
			36'b000000000000101010000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[30]=1'b1;
			end
			36'b000000000000010101000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[31]=1'b1;
			end
			36'b000000101010000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[32]=1'b1;
			end
			36'b000000010101000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[33]=1'b1;
			end
			36'b101010000000000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[34]=1'b1;
			end
			36'b010101000000000000000000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[35]=1'b1;
			end
			36'b000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			36'b100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_72_36_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [36-1:0] stored_data_edc = extended_hamming_code_72_36_f(i_stored_data);
wire [36-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [36-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_72_36_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_40_min_delay (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [40-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [40-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_80_40_f
//Compute 40 bits Error Detection Code from a 40 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 1208925819614629174706176 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[ 0]: x                                     x  (2 inputs)
//  syndrom[ 1]: x                                      x (2 inputs)
//  syndrom[ 2]:  x                                    x  (2 inputs)
//  syndrom[ 3]:  x                                     x (2 inputs)
//  syndrom[ 4]:   x                                 x    (2 inputs)
//  syndrom[ 5]:   x                                  x   (2 inputs)
//  syndrom[ 6]:    x                                x    (2 inputs)
//  syndrom[ 7]:    x                                 x   (2 inputs)
//  syndrom[ 8]:     x                             x      (2 inputs)
//  syndrom[ 9]:     x                              x     (2 inputs)
//  syndrom[10]:      x                            x      (2 inputs)
//  syndrom[11]:      x                             x     (2 inputs)
//  syndrom[12]:       x                         x        (2 inputs)
//  syndrom[13]:       x                          x       (2 inputs)
//  syndrom[14]:        x                        x        (2 inputs)
//  syndrom[15]:        x                         x       (2 inputs)
//  syndrom[16]:         x                     x          (2 inputs)
//  syndrom[17]:         x                      x         (2 inputs)
//  syndrom[18]:          x                    x          (2 inputs)
//  syndrom[19]:          x                     x         (2 inputs)
//  syndrom[20]:           x                 x            (2 inputs)
//  syndrom[21]:           x                  x           (2 inputs)
//  syndrom[22]:            x                x            (2 inputs)
//  syndrom[23]:            x                 x           (2 inputs)
//  syndrom[24]:             x             x              (2 inputs)
//  syndrom[25]:             x              x             (2 inputs)
//  syndrom[26]:              x            x              (2 inputs)
//  syndrom[27]:              x             x             (2 inputs)
//  syndrom[28]:               x         x                (2 inputs)
//  syndrom[29]:               x          x               (2 inputs)
//  syndrom[30]:                x        x                (2 inputs)
//  syndrom[31]:                x         x               (2 inputs)
//  syndrom[32]:                 x     x                  (2 inputs)
//  syndrom[33]:                 x      x                 (2 inputs)
//  syndrom[34]:                  x    x                  (2 inputs)
//  syndrom[35]:                  x     x                 (2 inputs)
//  syndrom[36]:                   x x                    (2 inputs)
//  syndrom[37]:                   x  x                   (2 inputs)
//  syndrom[38]:                    xx                    (2 inputs)
//  syndrom[39]:                    x x                   (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 32 33)
//  input bit 17 used  2 times (syndrom bits 34 35)
//  input bit 18 used  2 times (syndrom bits 36 37)
//  input bit 19 used  2 times (syndrom bits 38 39)
//  input bit 20 used  2 times (syndrom bits 36 38)
//  input bit 21 used  2 times (syndrom bits 37 39)
//  input bit 22 used  2 times (syndrom bits 32 34)
//  input bit 23 used  2 times (syndrom bits 33 35)
//  input bit 24 used  2 times (syndrom bits 28 30)
//  input bit 25 used  2 times (syndrom bits 29 31)
//  input bit 26 used  2 times (syndrom bits 24 26)
//  input bit 27 used  2 times (syndrom bits 25 27)
//  input bit 28 used  2 times (syndrom bits 20 22)
//  input bit 29 used  2 times (syndrom bits 21 23)
//  input bit 30 used  2 times (syndrom bits 16 18)
//  input bit 31 used  2 times (syndrom bits 17 19)
//  input bit 32 used  2 times (syndrom bits 12 14)
//  input bit 33 used  2 times (syndrom bits 13 15)
//  input bit 34 used  2 times (syndrom bits 8 10)
//  input bit 35 used  2 times (syndrom bits 9 11)
//  input bit 36 used  2 times (syndrom bits 4 6)
//  input bit 37 used  2 times (syndrom bits 5 7)
//  input bit 38 used  2 times (syndrom bits 0 2)
//  input bit 39 used  2 times (syndrom bits 1 3)
function [40-1:0] hamming_code_80_40_f;
    input [40-1:0] in;
    reg [40-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[38];//2 inputs
        syndrom[ 1] = in[ 0]^in[39];//2 inputs
        syndrom[ 2] = in[ 1]^in[38];//2 inputs
        syndrom[ 3] = in[ 1]^in[39];//2 inputs
        syndrom[ 4] = in[ 2]^in[36];//2 inputs
        syndrom[ 5] = in[ 2]^in[37];//2 inputs
        syndrom[ 6] = in[ 3]^in[36];//2 inputs
        syndrom[ 7] = in[ 3]^in[37];//2 inputs
        syndrom[ 8] = in[ 4]^in[34];//2 inputs
        syndrom[ 9] = in[ 4]^in[35];//2 inputs
        syndrom[10] = in[ 5]^in[34];//2 inputs
        syndrom[11] = in[ 5]^in[35];//2 inputs
        syndrom[12] = in[ 6]^in[32];//2 inputs
        syndrom[13] = in[ 6]^in[33];//2 inputs
        syndrom[14] = in[ 7]^in[32];//2 inputs
        syndrom[15] = in[ 7]^in[33];//2 inputs
        syndrom[16] = in[ 8]^in[30];//2 inputs
        syndrom[17] = in[ 8]^in[31];//2 inputs
        syndrom[18] = in[ 9]^in[30];//2 inputs
        syndrom[19] = in[ 9]^in[31];//2 inputs
        syndrom[20] = in[10]^in[28];//2 inputs
        syndrom[21] = in[10]^in[29];//2 inputs
        syndrom[22] = in[11]^in[28];//2 inputs
        syndrom[23] = in[11]^in[29];//2 inputs
        syndrom[24] = in[12]^in[26];//2 inputs
        syndrom[25] = in[12]^in[27];//2 inputs
        syndrom[26] = in[13]^in[26];//2 inputs
        syndrom[27] = in[13]^in[27];//2 inputs
        syndrom[28] = in[14]^in[24];//2 inputs
        syndrom[29] = in[14]^in[25];//2 inputs
        syndrom[30] = in[15]^in[24];//2 inputs
        syndrom[31] = in[15]^in[25];//2 inputs
        syndrom[32] = in[16]^in[22];//2 inputs
        syndrom[33] = in[16]^in[23];//2 inputs
        syndrom[34] = in[17]^in[22];//2 inputs
        syndrom[35] = in[17]^in[23];//2 inputs
        syndrom[36] = in[18]^in[20];//2 inputs
        syndrom[37] = in[18]^in[21];//2 inputs
        syndrom[38] = in[19]^in[20];//2 inputs
        syndrom[39] = in[19]^in[21];//2 inputs
        hamming_code_80_40_f = syndrom;
    end
endfunction
wire [40-1:0] stored_data_edc = hamming_code_80_40_f(i_stored_data);
wire [40-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_40_min_delay (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [40-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [40-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_80_40_f
//Compute 40 bits Error Detection Code from a 40 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 1208925819614629174706176 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[ 0]: x                        x  x            (3 inputs)
//  syndrom[ 1]: x                         xx             (3 inputs)
//  syndrom[ 2]: x                         xx             (3 inputs)
//  syndrom[ 3]:  x                      x    x           (3 inputs)
//  syndrom[ 4]:  x                       xx              (3 inputs)
//  syndrom[ 5]:  x                       x x             (3 inputs)
//  syndrom[ 6]:   x                    x      x          (3 inputs)
//  syndrom[ 7]:   x                     x   x            (3 inputs)
//  syndrom[ 8]:   x                     x   x            (3 inputs)
//  syndrom[ 9]:    x                  x        x         (3 inputs)
//  syndrom[10]:    x                   x     x           (3 inputs)
//  syndrom[11]:    x                   x     x           (3 inputs)
//  syndrom[12]:     x                x          x        (3 inputs)
//  syndrom[13]:     x                 x       x          (3 inputs)
//  syndrom[14]:     x                 x       x          (3 inputs)
//  syndrom[15]:      x              x            x       (3 inputs)
//  syndrom[16]:      x               x         x         (3 inputs)
//  syndrom[17]:      x               x         x         (3 inputs)
//  syndrom[18]:       x            x              x      (3 inputs)
//  syndrom[19]:       x             x           x        (3 inputs)
//  syndrom[20]:       x             x           x        (3 inputs)
//  syndrom[21]:        x          x                x     (3 inputs)
//  syndrom[22]:        x           x             x       (3 inputs)
//  syndrom[23]:        x           x             x       (3 inputs)
//  syndrom[24]:         x        x                  x    (3 inputs)
//  syndrom[25]:         x         x               x      (3 inputs)
//  syndrom[26]:         x         x               x      (3 inputs)
//  syndrom[27]:          x      x                    x   (3 inputs)
//  syndrom[28]:          x       x                 x     (3 inputs)
//  syndrom[29]:          x       x                 x     (3 inputs)
//  syndrom[30]:           x    x                      x  (3 inputs)
//  syndrom[31]:           x     x                   x    (3 inputs)
//  syndrom[32]:           x     x                   x    (3 inputs)
//  syndrom[33]:            x  x                        x (3 inputs)
//  syndrom[34]:            x   x                     x   (3 inputs)
//  syndrom[35]:            x   x                     x   (3 inputs)
//  syndrom[36]:             xx                         x (3 inputs)
//  syndrom[37]:             xx                         x (3 inputs)
//  syndrom[38]:             x x                       x  (3 inputs)
//  syndrom[39]:              xx                       x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 36 37 39)
//  input bit 14 used  3 times (syndrom bits 33 38 39)
//  input bit 15 used  3 times (syndrom bits 30 34 35)
//  input bit 16 used  3 times (syndrom bits 27 31 32)
//  input bit 17 used  3 times (syndrom bits 24 28 29)
//  input bit 18 used  3 times (syndrom bits 21 25 26)
//  input bit 19 used  3 times (syndrom bits 18 22 23)
//  input bit 20 used  3 times (syndrom bits 15 19 20)
//  input bit 21 used  3 times (syndrom bits 12 16 17)
//  input bit 22 used  3 times (syndrom bits 9 13 14)
//  input bit 23 used  3 times (syndrom bits 6 10 11)
//  input bit 24 used  3 times (syndrom bits 3 7 8)
//  input bit 25 used  3 times (syndrom bits 0 4 5)
//  input bit 26 used  3 times (syndrom bits 1 2 4)
//  input bit 27 used  3 times (syndrom bits 1 2 5)
//  input bit 28 used  3 times (syndrom bits 0 7 8)
//  input bit 29 used  3 times (syndrom bits 3 10 11)
//  input bit 30 used  3 times (syndrom bits 6 13 14)
//  input bit 31 used  3 times (syndrom bits 9 16 17)
//  input bit 32 used  3 times (syndrom bits 12 19 20)
//  input bit 33 used  3 times (syndrom bits 15 22 23)
//  input bit 34 used  3 times (syndrom bits 18 25 26)
//  input bit 35 used  3 times (syndrom bits 21 28 29)
//  input bit 36 used  3 times (syndrom bits 24 31 32)
//  input bit 37 used  3 times (syndrom bits 27 34 35)
//  input bit 38 used  3 times (syndrom bits 30 38 39)
//  input bit 39 used  3 times (syndrom bits 33 36 37)
function [40-1:0] extended_hamming_code_80_40_f;
    input [40-1:0] in;
    reg [40-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[25]^in[28];//3 inputs
        syndrom[ 1] = in[ 0]^in[26]^in[27];//3 inputs
        syndrom[ 2] = in[ 0]^in[26]^in[27];//3 inputs
        syndrom[ 3] = in[ 1]^in[24]^in[29];//3 inputs
        syndrom[ 4] = in[ 1]^in[25]^in[26];//3 inputs
        syndrom[ 5] = in[ 1]^in[25]^in[27];//3 inputs
        syndrom[ 6] = in[ 2]^in[23]^in[30];//3 inputs
        syndrom[ 7] = in[ 2]^in[24]^in[28];//3 inputs
        syndrom[ 8] = in[ 2]^in[24]^in[28];//3 inputs
        syndrom[ 9] = in[ 3]^in[22]^in[31];//3 inputs
        syndrom[10] = in[ 3]^in[23]^in[29];//3 inputs
        syndrom[11] = in[ 3]^in[23]^in[29];//3 inputs
        syndrom[12] = in[ 4]^in[21]^in[32];//3 inputs
        syndrom[13] = in[ 4]^in[22]^in[30];//3 inputs
        syndrom[14] = in[ 4]^in[22]^in[30];//3 inputs
        syndrom[15] = in[ 5]^in[20]^in[33];//3 inputs
        syndrom[16] = in[ 5]^in[21]^in[31];//3 inputs
        syndrom[17] = in[ 5]^in[21]^in[31];//3 inputs
        syndrom[18] = in[ 6]^in[19]^in[34];//3 inputs
        syndrom[19] = in[ 6]^in[20]^in[32];//3 inputs
        syndrom[20] = in[ 6]^in[20]^in[32];//3 inputs
        syndrom[21] = in[ 7]^in[18]^in[35];//3 inputs
        syndrom[22] = in[ 7]^in[19]^in[33];//3 inputs
        syndrom[23] = in[ 7]^in[19]^in[33];//3 inputs
        syndrom[24] = in[ 8]^in[17]^in[36];//3 inputs
        syndrom[25] = in[ 8]^in[18]^in[34];//3 inputs
        syndrom[26] = in[ 8]^in[18]^in[34];//3 inputs
        syndrom[27] = in[ 9]^in[16]^in[37];//3 inputs
        syndrom[28] = in[ 9]^in[17]^in[35];//3 inputs
        syndrom[29] = in[ 9]^in[17]^in[35];//3 inputs
        syndrom[30] = in[10]^in[15]^in[38];//3 inputs
        syndrom[31] = in[10]^in[16]^in[36];//3 inputs
        syndrom[32] = in[10]^in[16]^in[36];//3 inputs
        syndrom[33] = in[11]^in[14]^in[39];//3 inputs
        syndrom[34] = in[11]^in[15]^in[37];//3 inputs
        syndrom[35] = in[11]^in[15]^in[37];//3 inputs
        syndrom[36] = in[12]^in[13]^in[39];//3 inputs
        syndrom[37] = in[12]^in[13]^in[39];//3 inputs
        syndrom[38] = in[12]^in[14]^in[38];//3 inputs
        syndrom[39] = in[13]^in[14]^in[38];//3 inputs
        extended_hamming_code_80_40_f = syndrom;
    end
endfunction
wire [40-1:0] stored_data_edc = extended_hamming_code_80_40_f(i_stored_data);
wire [40-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_40_min_delay (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [40-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [40-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [40-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_80_40_f
//Compute 40 bits Error Detection Code from a 40 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 1208925819614629174706176 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[ 0]: x                        x  x            (3 inputs)
//  syndrom[ 1]: x                         xx             (3 inputs)
//  syndrom[ 2]: x                         xx             (3 inputs)
//  syndrom[ 3]:  x                      x    x           (3 inputs)
//  syndrom[ 4]:  x                       xx              (3 inputs)
//  syndrom[ 5]:  x                       x x             (3 inputs)
//  syndrom[ 6]:   x                    x      x          (3 inputs)
//  syndrom[ 7]:   x                     x   x            (3 inputs)
//  syndrom[ 8]:   x                     x   x            (3 inputs)
//  syndrom[ 9]:    x                  x        x         (3 inputs)
//  syndrom[10]:    x                   x     x           (3 inputs)
//  syndrom[11]:    x                   x     x           (3 inputs)
//  syndrom[12]:     x                x          x        (3 inputs)
//  syndrom[13]:     x                 x       x          (3 inputs)
//  syndrom[14]:     x                 x       x          (3 inputs)
//  syndrom[15]:      x              x            x       (3 inputs)
//  syndrom[16]:      x               x         x         (3 inputs)
//  syndrom[17]:      x               x         x         (3 inputs)
//  syndrom[18]:       x            x              x      (3 inputs)
//  syndrom[19]:       x             x           x        (3 inputs)
//  syndrom[20]:       x             x           x        (3 inputs)
//  syndrom[21]:        x          x                x     (3 inputs)
//  syndrom[22]:        x           x             x       (3 inputs)
//  syndrom[23]:        x           x             x       (3 inputs)
//  syndrom[24]:         x        x                  x    (3 inputs)
//  syndrom[25]:         x         x               x      (3 inputs)
//  syndrom[26]:         x         x               x      (3 inputs)
//  syndrom[27]:          x      x                    x   (3 inputs)
//  syndrom[28]:          x       x                 x     (3 inputs)
//  syndrom[29]:          x       x                 x     (3 inputs)
//  syndrom[30]:           x    x                      x  (3 inputs)
//  syndrom[31]:           x     x                   x    (3 inputs)
//  syndrom[32]:           x     x                   x    (3 inputs)
//  syndrom[33]:            x  x                        x (3 inputs)
//  syndrom[34]:            x   x                     x   (3 inputs)
//  syndrom[35]:            x   x                     x   (3 inputs)
//  syndrom[36]:             xx                         x (3 inputs)
//  syndrom[37]:             xx                         x (3 inputs)
//  syndrom[38]:             x x                       x  (3 inputs)
//  syndrom[39]:              xx                       x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 36 37 39)
//  input bit 14 used  3 times (syndrom bits 33 38 39)
//  input bit 15 used  3 times (syndrom bits 30 34 35)
//  input bit 16 used  3 times (syndrom bits 27 31 32)
//  input bit 17 used  3 times (syndrom bits 24 28 29)
//  input bit 18 used  3 times (syndrom bits 21 25 26)
//  input bit 19 used  3 times (syndrom bits 18 22 23)
//  input bit 20 used  3 times (syndrom bits 15 19 20)
//  input bit 21 used  3 times (syndrom bits 12 16 17)
//  input bit 22 used  3 times (syndrom bits 9 13 14)
//  input bit 23 used  3 times (syndrom bits 6 10 11)
//  input bit 24 used  3 times (syndrom bits 3 7 8)
//  input bit 25 used  3 times (syndrom bits 0 4 5)
//  input bit 26 used  3 times (syndrom bits 1 2 4)
//  input bit 27 used  3 times (syndrom bits 1 2 5)
//  input bit 28 used  3 times (syndrom bits 0 7 8)
//  input bit 29 used  3 times (syndrom bits 3 10 11)
//  input bit 30 used  3 times (syndrom bits 6 13 14)
//  input bit 31 used  3 times (syndrom bits 9 16 17)
//  input bit 32 used  3 times (syndrom bits 12 19 20)
//  input bit 33 used  3 times (syndrom bits 15 22 23)
//  input bit 34 used  3 times (syndrom bits 18 25 26)
//  input bit 35 used  3 times (syndrom bits 21 28 29)
//  input bit 36 used  3 times (syndrom bits 24 31 32)
//  input bit 37 used  3 times (syndrom bits 27 34 35)
//  input bit 38 used  3 times (syndrom bits 30 38 39)
//  input bit 39 used  3 times (syndrom bits 33 36 37)
function [40-1:0] extended_hamming_code_80_40_f;
    input [40-1:0] in;
    reg [40-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[25]^in[28];//3 inputs
        syndrom[ 1] = in[ 0]^in[26]^in[27];//3 inputs
        syndrom[ 2] = in[ 0]^in[26]^in[27];//3 inputs
        syndrom[ 3] = in[ 1]^in[24]^in[29];//3 inputs
        syndrom[ 4] = in[ 1]^in[25]^in[26];//3 inputs
        syndrom[ 5] = in[ 1]^in[25]^in[27];//3 inputs
        syndrom[ 6] = in[ 2]^in[23]^in[30];//3 inputs
        syndrom[ 7] = in[ 2]^in[24]^in[28];//3 inputs
        syndrom[ 8] = in[ 2]^in[24]^in[28];//3 inputs
        syndrom[ 9] = in[ 3]^in[22]^in[31];//3 inputs
        syndrom[10] = in[ 3]^in[23]^in[29];//3 inputs
        syndrom[11] = in[ 3]^in[23]^in[29];//3 inputs
        syndrom[12] = in[ 4]^in[21]^in[32];//3 inputs
        syndrom[13] = in[ 4]^in[22]^in[30];//3 inputs
        syndrom[14] = in[ 4]^in[22]^in[30];//3 inputs
        syndrom[15] = in[ 5]^in[20]^in[33];//3 inputs
        syndrom[16] = in[ 5]^in[21]^in[31];//3 inputs
        syndrom[17] = in[ 5]^in[21]^in[31];//3 inputs
        syndrom[18] = in[ 6]^in[19]^in[34];//3 inputs
        syndrom[19] = in[ 6]^in[20]^in[32];//3 inputs
        syndrom[20] = in[ 6]^in[20]^in[32];//3 inputs
        syndrom[21] = in[ 7]^in[18]^in[35];//3 inputs
        syndrom[22] = in[ 7]^in[19]^in[33];//3 inputs
        syndrom[23] = in[ 7]^in[19]^in[33];//3 inputs
        syndrom[24] = in[ 8]^in[17]^in[36];//3 inputs
        syndrom[25] = in[ 8]^in[18]^in[34];//3 inputs
        syndrom[26] = in[ 8]^in[18]^in[34];//3 inputs
        syndrom[27] = in[ 9]^in[16]^in[37];//3 inputs
        syndrom[28] = in[ 9]^in[17]^in[35];//3 inputs
        syndrom[29] = in[ 9]^in[17]^in[35];//3 inputs
        syndrom[30] = in[10]^in[15]^in[38];//3 inputs
        syndrom[31] = in[10]^in[16]^in[36];//3 inputs
        syndrom[32] = in[10]^in[16]^in[36];//3 inputs
        syndrom[33] = in[11]^in[14]^in[39];//3 inputs
        syndrom[34] = in[11]^in[15]^in[37];//3 inputs
        syndrom[35] = in[11]^in[15]^in[37];//3 inputs
        syndrom[36] = in[12]^in[13]^in[39];//3 inputs
        syndrom[37] = in[12]^in[13]^in[39];//3 inputs
        syndrom[38] = in[12]^in[14]^in[38];//3 inputs
        syndrom[39] = in[13]^in[14]^in[38];//3 inputs
        extended_hamming_code_80_40_f = syndrom;
    end
endfunction
function [2+40-1:0] extended_hamming_code_80_40_f_correction_pattern_f;
    input [40-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [40-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {40{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			40'b0000000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {40{1'b0}};
			end	
			40'b0000000000000000000000000000000000000111: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 0]=1'b1;
			end
			40'b0000000000000000000000000000000000111000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 1]=1'b1;
			end
			40'b0000000000000000000000000000000111000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 2]=1'b1;
			end
			40'b0000000000000000000000000000111000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 3]=1'b1;
			end
			40'b0000000000000000000000000111000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 4]=1'b1;
			end
			40'b0000000000000000000000111000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 5]=1'b1;
			end
			40'b0000000000000000000111000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 6]=1'b1;
			end
			40'b0000000000000000111000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 7]=1'b1;
			end
			40'b0000000000000111000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 8]=1'b1;
			end
			40'b0000000000111000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 9]=1'b1;
			end
			40'b0000000111000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[10]=1'b1;
			end
			40'b0000111000000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[11]=1'b1;
			end
			40'b0111000000000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[12]=1'b1;
			end
			40'b1011000000000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[13]=1'b1;
			end
			40'b1100001000000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[14]=1'b1;
			end
			40'b0000110001000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[15]=1'b1;
			end
			40'b0000000110001000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[16]=1'b1;
			end
			40'b0000000000110001000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[17]=1'b1;
			end
			40'b0000000000000110001000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[18]=1'b1;
			end
			40'b0000000000000000110001000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[19]=1'b1;
			end
			40'b0000000000000000000110001000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[20]=1'b1;
			end
			40'b0000000000000000000000110001000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[21]=1'b1;
			end
			40'b0000000000000000000000000110001000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[22]=1'b1;
			end
			40'b0000000000000000000000000000110001000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[23]=1'b1;
			end
			40'b0000000000000000000000000000000110001000: begin
				correction_pattern = {40{1'b0}};correction_pattern[24]=1'b1;
			end
			40'b0000000000000000000000000000000000110001: begin
				correction_pattern = {40{1'b0}};correction_pattern[25]=1'b1;
			end
			40'b0000000000000000000000000000000000010110: begin
				correction_pattern = {40{1'b0}};correction_pattern[26]=1'b1;
			end
			40'b0000000000000000000000000000000000100110: begin
				correction_pattern = {40{1'b0}};correction_pattern[27]=1'b1;
			end
			40'b0000000000000000000000000000000110000001: begin
				correction_pattern = {40{1'b0}};correction_pattern[28]=1'b1;
			end
			40'b0000000000000000000000000000110000001000: begin
				correction_pattern = {40{1'b0}};correction_pattern[29]=1'b1;
			end
			40'b0000000000000000000000000110000001000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[30]=1'b1;
			end
			40'b0000000000000000000000110000001000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[31]=1'b1;
			end
			40'b0000000000000000000110000001000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[32]=1'b1;
			end
			40'b0000000000000000110000001000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[33]=1'b1;
			end
			40'b0000000000000110000001000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[34]=1'b1;
			end
			40'b0000000000110000001000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[35]=1'b1;
			end
			40'b0000000110000001000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[36]=1'b1;
			end
			40'b0000110000001000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[37]=1'b1;
			end
			40'b1100000001000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[38]=1'b1;
			end
			40'b0011001000000000000000000000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[39]=1'b1;
			end
			40'b0000000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0000100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0001000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0010000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b0100000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			40'b1000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_80_40_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [40-1:0] stored_data_edc = extended_hamming_code_80_40_f(i_stored_data);
wire [40-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [40-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_80_40_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_48_min_delay (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [48-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [48-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_96_48_f
//Compute 48 bits Error Detection Code from a 48 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 79228162514264337593543950336 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[ 0]: x                                             x  (2 inputs)
//  syndrom[ 1]: x                                              x (2 inputs)
//  syndrom[ 2]:  x                                            x  (2 inputs)
//  syndrom[ 3]:  x                                             x (2 inputs)
//  syndrom[ 4]:   x                                         x    (2 inputs)
//  syndrom[ 5]:   x                                          x   (2 inputs)
//  syndrom[ 6]:    x                                        x    (2 inputs)
//  syndrom[ 7]:    x                                         x   (2 inputs)
//  syndrom[ 8]:     x                                     x      (2 inputs)
//  syndrom[ 9]:     x                                      x     (2 inputs)
//  syndrom[10]:      x                                    x      (2 inputs)
//  syndrom[11]:      x                                     x     (2 inputs)
//  syndrom[12]:       x                                 x        (2 inputs)
//  syndrom[13]:       x                                  x       (2 inputs)
//  syndrom[14]:        x                                x        (2 inputs)
//  syndrom[15]:        x                                 x       (2 inputs)
//  syndrom[16]:         x                             x          (2 inputs)
//  syndrom[17]:         x                              x         (2 inputs)
//  syndrom[18]:          x                            x          (2 inputs)
//  syndrom[19]:          x                             x         (2 inputs)
//  syndrom[20]:           x                         x            (2 inputs)
//  syndrom[21]:           x                          x           (2 inputs)
//  syndrom[22]:            x                        x            (2 inputs)
//  syndrom[23]:            x                         x           (2 inputs)
//  syndrom[24]:             x                     x              (2 inputs)
//  syndrom[25]:             x                      x             (2 inputs)
//  syndrom[26]:              x                    x              (2 inputs)
//  syndrom[27]:              x                     x             (2 inputs)
//  syndrom[28]:               x                 x                (2 inputs)
//  syndrom[29]:               x                  x               (2 inputs)
//  syndrom[30]:                x                x                (2 inputs)
//  syndrom[31]:                x                 x               (2 inputs)
//  syndrom[32]:                 x             x                  (2 inputs)
//  syndrom[33]:                 x              x                 (2 inputs)
//  syndrom[34]:                  x            x                  (2 inputs)
//  syndrom[35]:                  x             x                 (2 inputs)
//  syndrom[36]:                   x         x                    (2 inputs)
//  syndrom[37]:                   x          x                   (2 inputs)
//  syndrom[38]:                    x        x                    (2 inputs)
//  syndrom[39]:                    x         x                   (2 inputs)
//  syndrom[40]:                     x     x                      (2 inputs)
//  syndrom[41]:                     x      x                     (2 inputs)
//  syndrom[42]:                      x    x                      (2 inputs)
//  syndrom[43]:                      x     x                     (2 inputs)
//  syndrom[44]:                       x x                        (2 inputs)
//  syndrom[45]:                       x  x                       (2 inputs)
//  syndrom[46]:                        xx                        (2 inputs)
//  syndrom[47]:                        x x                       (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 32 33)
//  input bit 17 used  2 times (syndrom bits 34 35)
//  input bit 18 used  2 times (syndrom bits 36 37)
//  input bit 19 used  2 times (syndrom bits 38 39)
//  input bit 20 used  2 times (syndrom bits 40 41)
//  input bit 21 used  2 times (syndrom bits 42 43)
//  input bit 22 used  2 times (syndrom bits 44 45)
//  input bit 23 used  2 times (syndrom bits 46 47)
//  input bit 24 used  2 times (syndrom bits 44 46)
//  input bit 25 used  2 times (syndrom bits 45 47)
//  input bit 26 used  2 times (syndrom bits 40 42)
//  input bit 27 used  2 times (syndrom bits 41 43)
//  input bit 28 used  2 times (syndrom bits 36 38)
//  input bit 29 used  2 times (syndrom bits 37 39)
//  input bit 30 used  2 times (syndrom bits 32 34)
//  input bit 31 used  2 times (syndrom bits 33 35)
//  input bit 32 used  2 times (syndrom bits 28 30)
//  input bit 33 used  2 times (syndrom bits 29 31)
//  input bit 34 used  2 times (syndrom bits 24 26)
//  input bit 35 used  2 times (syndrom bits 25 27)
//  input bit 36 used  2 times (syndrom bits 20 22)
//  input bit 37 used  2 times (syndrom bits 21 23)
//  input bit 38 used  2 times (syndrom bits 16 18)
//  input bit 39 used  2 times (syndrom bits 17 19)
//  input bit 40 used  2 times (syndrom bits 12 14)
//  input bit 41 used  2 times (syndrom bits 13 15)
//  input bit 42 used  2 times (syndrom bits 8 10)
//  input bit 43 used  2 times (syndrom bits 9 11)
//  input bit 44 used  2 times (syndrom bits 4 6)
//  input bit 45 used  2 times (syndrom bits 5 7)
//  input bit 46 used  2 times (syndrom bits 0 2)
//  input bit 47 used  2 times (syndrom bits 1 3)
function [48-1:0] hamming_code_96_48_f;
    input [48-1:0] in;
    reg [48-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[46];//2 inputs
        syndrom[ 1] = in[ 0]^in[47];//2 inputs
        syndrom[ 2] = in[ 1]^in[46];//2 inputs
        syndrom[ 3] = in[ 1]^in[47];//2 inputs
        syndrom[ 4] = in[ 2]^in[44];//2 inputs
        syndrom[ 5] = in[ 2]^in[45];//2 inputs
        syndrom[ 6] = in[ 3]^in[44];//2 inputs
        syndrom[ 7] = in[ 3]^in[45];//2 inputs
        syndrom[ 8] = in[ 4]^in[42];//2 inputs
        syndrom[ 9] = in[ 4]^in[43];//2 inputs
        syndrom[10] = in[ 5]^in[42];//2 inputs
        syndrom[11] = in[ 5]^in[43];//2 inputs
        syndrom[12] = in[ 6]^in[40];//2 inputs
        syndrom[13] = in[ 6]^in[41];//2 inputs
        syndrom[14] = in[ 7]^in[40];//2 inputs
        syndrom[15] = in[ 7]^in[41];//2 inputs
        syndrom[16] = in[ 8]^in[38];//2 inputs
        syndrom[17] = in[ 8]^in[39];//2 inputs
        syndrom[18] = in[ 9]^in[38];//2 inputs
        syndrom[19] = in[ 9]^in[39];//2 inputs
        syndrom[20] = in[10]^in[36];//2 inputs
        syndrom[21] = in[10]^in[37];//2 inputs
        syndrom[22] = in[11]^in[36];//2 inputs
        syndrom[23] = in[11]^in[37];//2 inputs
        syndrom[24] = in[12]^in[34];//2 inputs
        syndrom[25] = in[12]^in[35];//2 inputs
        syndrom[26] = in[13]^in[34];//2 inputs
        syndrom[27] = in[13]^in[35];//2 inputs
        syndrom[28] = in[14]^in[32];//2 inputs
        syndrom[29] = in[14]^in[33];//2 inputs
        syndrom[30] = in[15]^in[32];//2 inputs
        syndrom[31] = in[15]^in[33];//2 inputs
        syndrom[32] = in[16]^in[30];//2 inputs
        syndrom[33] = in[16]^in[31];//2 inputs
        syndrom[34] = in[17]^in[30];//2 inputs
        syndrom[35] = in[17]^in[31];//2 inputs
        syndrom[36] = in[18]^in[28];//2 inputs
        syndrom[37] = in[18]^in[29];//2 inputs
        syndrom[38] = in[19]^in[28];//2 inputs
        syndrom[39] = in[19]^in[29];//2 inputs
        syndrom[40] = in[20]^in[26];//2 inputs
        syndrom[41] = in[20]^in[27];//2 inputs
        syndrom[42] = in[21]^in[26];//2 inputs
        syndrom[43] = in[21]^in[27];//2 inputs
        syndrom[44] = in[22]^in[24];//2 inputs
        syndrom[45] = in[22]^in[25];//2 inputs
        syndrom[46] = in[23]^in[24];//2 inputs
        syndrom[47] = in[23]^in[25];//2 inputs
        hamming_code_96_48_f = syndrom;
    end
endfunction
wire [48-1:0] stored_data_edc = hamming_code_96_48_f(i_stored_data);
wire [48-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_48_min_delay (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [48-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [48-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_96_48_f
//Compute 48 bits Error Detection Code from a 48 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 79228162514264337593543950336 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[ 0]: x                             x  x               (3 inputs)
//  syndrom[ 1]: x                              xx                (3 inputs)
//  syndrom[ 2]: x                              x x               (3 inputs)
//  syndrom[ 3]:  x                            x x                (3 inputs)
//  syndrom[ 4]:  x                            x  x               (3 inputs)
//  syndrom[ 5]:  x                             xx                (3 inputs)
//  syndrom[ 6]:   x                         x      x             (3 inputs)
//  syndrom[ 7]:   x                          x    x              (3 inputs)
//  syndrom[ 8]:   x                          x     x             (3 inputs)
//  syndrom[ 9]:    x                        x     x              (3 inputs)
//  syndrom[10]:    x                        x      x             (3 inputs)
//  syndrom[11]:    x                         x    x              (3 inputs)
//  syndrom[12]:     x                     x          x           (3 inputs)
//  syndrom[13]:     x                      x        x            (3 inputs)
//  syndrom[14]:     x                      x         x           (3 inputs)
//  syndrom[15]:      x                    x         x            (3 inputs)
//  syndrom[16]:      x                    x          x           (3 inputs)
//  syndrom[17]:      x                     x        x            (3 inputs)
//  syndrom[18]:       x                 x              x         (3 inputs)
//  syndrom[19]:       x                  x            x          (3 inputs)
//  syndrom[20]:       x                  x             x         (3 inputs)
//  syndrom[21]:        x                x             x          (3 inputs)
//  syndrom[22]:        x                x              x         (3 inputs)
//  syndrom[23]:        x                 x            x          (3 inputs)
//  syndrom[24]:         x             x                  x       (3 inputs)
//  syndrom[25]:         x              x                x        (3 inputs)
//  syndrom[26]:         x              x                 x       (3 inputs)
//  syndrom[27]:          x            x                 x        (3 inputs)
//  syndrom[28]:          x            x                  x       (3 inputs)
//  syndrom[29]:          x             x                x        (3 inputs)
//  syndrom[30]:           x         x                      x     (3 inputs)
//  syndrom[31]:           x          x                    x      (3 inputs)
//  syndrom[32]:           x          x                     x     (3 inputs)
//  syndrom[33]:            x        x                     x      (3 inputs)
//  syndrom[34]:            x        x                      x     (3 inputs)
//  syndrom[35]:            x         x                    x      (3 inputs)
//  syndrom[36]:             x     x                          x   (3 inputs)
//  syndrom[37]:             x      x                        x    (3 inputs)
//  syndrom[38]:             x      x                         x   (3 inputs)
//  syndrom[39]:              x    x                         x    (3 inputs)
//  syndrom[40]:              x    x                          x   (3 inputs)
//  syndrom[41]:              x     x                        x    (3 inputs)
//  syndrom[42]:               x x                              x (3 inputs)
//  syndrom[43]:               x  x                            x  (3 inputs)
//  syndrom[44]:               x  x                             x (3 inputs)
//  syndrom[45]:                xx                             x  (3 inputs)
//  syndrom[46]:                xx                              x (3 inputs)
//  syndrom[47]:                x x                            x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 42 45 46)
//  input bit 17 used  3 times (syndrom bits 43 44 47)
//  input bit 18 used  3 times (syndrom bits 36 39 40)
//  input bit 19 used  3 times (syndrom bits 37 38 41)
//  input bit 20 used  3 times (syndrom bits 30 33 34)
//  input bit 21 used  3 times (syndrom bits 31 32 35)
//  input bit 22 used  3 times (syndrom bits 24 27 28)
//  input bit 23 used  3 times (syndrom bits 25 26 29)
//  input bit 24 used  3 times (syndrom bits 18 21 22)
//  input bit 25 used  3 times (syndrom bits 19 20 23)
//  input bit 26 used  3 times (syndrom bits 12 15 16)
//  input bit 27 used  3 times (syndrom bits 13 14 17)
//  input bit 28 used  3 times (syndrom bits 6 9 10)
//  input bit 29 used  3 times (syndrom bits 7 8 11)
//  input bit 30 used  3 times (syndrom bits 0 3 4)
//  input bit 31 used  3 times (syndrom bits 1 2 5)
//  input bit 32 used  3 times (syndrom bits 1 3 5)
//  input bit 33 used  3 times (syndrom bits 0 2 4)
//  input bit 34 used  3 times (syndrom bits 7 9 11)
//  input bit 35 used  3 times (syndrom bits 6 8 10)
//  input bit 36 used  3 times (syndrom bits 13 15 17)
//  input bit 37 used  3 times (syndrom bits 12 14 16)
//  input bit 38 used  3 times (syndrom bits 19 21 23)
//  input bit 39 used  3 times (syndrom bits 18 20 22)
//  input bit 40 used  3 times (syndrom bits 25 27 29)
//  input bit 41 used  3 times (syndrom bits 24 26 28)
//  input bit 42 used  3 times (syndrom bits 31 33 35)
//  input bit 43 used  3 times (syndrom bits 30 32 34)
//  input bit 44 used  3 times (syndrom bits 37 39 41)
//  input bit 45 used  3 times (syndrom bits 36 38 40)
//  input bit 46 used  3 times (syndrom bits 43 45 47)
//  input bit 47 used  3 times (syndrom bits 42 44 46)
function [48-1:0] extended_hamming_code_96_48_f;
    input [48-1:0] in;
    reg [48-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[30]^in[33];//3 inputs
        syndrom[ 1] = in[ 0]^in[31]^in[32];//3 inputs
        syndrom[ 2] = in[ 0]^in[31]^in[33];//3 inputs
        syndrom[ 3] = in[ 1]^in[30]^in[32];//3 inputs
        syndrom[ 4] = in[ 1]^in[30]^in[33];//3 inputs
        syndrom[ 5] = in[ 1]^in[31]^in[32];//3 inputs
        syndrom[ 6] = in[ 2]^in[28]^in[35];//3 inputs
        syndrom[ 7] = in[ 2]^in[29]^in[34];//3 inputs
        syndrom[ 8] = in[ 2]^in[29]^in[35];//3 inputs
        syndrom[ 9] = in[ 3]^in[28]^in[34];//3 inputs
        syndrom[10] = in[ 3]^in[28]^in[35];//3 inputs
        syndrom[11] = in[ 3]^in[29]^in[34];//3 inputs
        syndrom[12] = in[ 4]^in[26]^in[37];//3 inputs
        syndrom[13] = in[ 4]^in[27]^in[36];//3 inputs
        syndrom[14] = in[ 4]^in[27]^in[37];//3 inputs
        syndrom[15] = in[ 5]^in[26]^in[36];//3 inputs
        syndrom[16] = in[ 5]^in[26]^in[37];//3 inputs
        syndrom[17] = in[ 5]^in[27]^in[36];//3 inputs
        syndrom[18] = in[ 6]^in[24]^in[39];//3 inputs
        syndrom[19] = in[ 6]^in[25]^in[38];//3 inputs
        syndrom[20] = in[ 6]^in[25]^in[39];//3 inputs
        syndrom[21] = in[ 7]^in[24]^in[38];//3 inputs
        syndrom[22] = in[ 7]^in[24]^in[39];//3 inputs
        syndrom[23] = in[ 7]^in[25]^in[38];//3 inputs
        syndrom[24] = in[ 8]^in[22]^in[41];//3 inputs
        syndrom[25] = in[ 8]^in[23]^in[40];//3 inputs
        syndrom[26] = in[ 8]^in[23]^in[41];//3 inputs
        syndrom[27] = in[ 9]^in[22]^in[40];//3 inputs
        syndrom[28] = in[ 9]^in[22]^in[41];//3 inputs
        syndrom[29] = in[ 9]^in[23]^in[40];//3 inputs
        syndrom[30] = in[10]^in[20]^in[43];//3 inputs
        syndrom[31] = in[10]^in[21]^in[42];//3 inputs
        syndrom[32] = in[10]^in[21]^in[43];//3 inputs
        syndrom[33] = in[11]^in[20]^in[42];//3 inputs
        syndrom[34] = in[11]^in[20]^in[43];//3 inputs
        syndrom[35] = in[11]^in[21]^in[42];//3 inputs
        syndrom[36] = in[12]^in[18]^in[45];//3 inputs
        syndrom[37] = in[12]^in[19]^in[44];//3 inputs
        syndrom[38] = in[12]^in[19]^in[45];//3 inputs
        syndrom[39] = in[13]^in[18]^in[44];//3 inputs
        syndrom[40] = in[13]^in[18]^in[45];//3 inputs
        syndrom[41] = in[13]^in[19]^in[44];//3 inputs
        syndrom[42] = in[14]^in[16]^in[47];//3 inputs
        syndrom[43] = in[14]^in[17]^in[46];//3 inputs
        syndrom[44] = in[14]^in[17]^in[47];//3 inputs
        syndrom[45] = in[15]^in[16]^in[46];//3 inputs
        syndrom[46] = in[15]^in[16]^in[47];//3 inputs
        syndrom[47] = in[15]^in[17]^in[46];//3 inputs
        extended_hamming_code_96_48_f = syndrom;
    end
endfunction
wire [48-1:0] stored_data_edc = extended_hamming_code_96_48_f(i_stored_data);
wire [48-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_48_min_delay (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [48-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [48-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [48-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_96_48_f
//Compute 48 bits Error Detection Code from a 48 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 79228162514264337593543950336 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[ 0]: x                             x  x               (3 inputs)
//  syndrom[ 1]: x                              xx                (3 inputs)
//  syndrom[ 2]: x                              x x               (3 inputs)
//  syndrom[ 3]:  x                            x x                (3 inputs)
//  syndrom[ 4]:  x                            x  x               (3 inputs)
//  syndrom[ 5]:  x                             xx                (3 inputs)
//  syndrom[ 6]:   x                         x      x             (3 inputs)
//  syndrom[ 7]:   x                          x    x              (3 inputs)
//  syndrom[ 8]:   x                          x     x             (3 inputs)
//  syndrom[ 9]:    x                        x     x              (3 inputs)
//  syndrom[10]:    x                        x      x             (3 inputs)
//  syndrom[11]:    x                         x    x              (3 inputs)
//  syndrom[12]:     x                     x          x           (3 inputs)
//  syndrom[13]:     x                      x        x            (3 inputs)
//  syndrom[14]:     x                      x         x           (3 inputs)
//  syndrom[15]:      x                    x         x            (3 inputs)
//  syndrom[16]:      x                    x          x           (3 inputs)
//  syndrom[17]:      x                     x        x            (3 inputs)
//  syndrom[18]:       x                 x              x         (3 inputs)
//  syndrom[19]:       x                  x            x          (3 inputs)
//  syndrom[20]:       x                  x             x         (3 inputs)
//  syndrom[21]:        x                x             x          (3 inputs)
//  syndrom[22]:        x                x              x         (3 inputs)
//  syndrom[23]:        x                 x            x          (3 inputs)
//  syndrom[24]:         x             x                  x       (3 inputs)
//  syndrom[25]:         x              x                x        (3 inputs)
//  syndrom[26]:         x              x                 x       (3 inputs)
//  syndrom[27]:          x            x                 x        (3 inputs)
//  syndrom[28]:          x            x                  x       (3 inputs)
//  syndrom[29]:          x             x                x        (3 inputs)
//  syndrom[30]:           x         x                      x     (3 inputs)
//  syndrom[31]:           x          x                    x      (3 inputs)
//  syndrom[32]:           x          x                     x     (3 inputs)
//  syndrom[33]:            x        x                     x      (3 inputs)
//  syndrom[34]:            x        x                      x     (3 inputs)
//  syndrom[35]:            x         x                    x      (3 inputs)
//  syndrom[36]:             x     x                          x   (3 inputs)
//  syndrom[37]:             x      x                        x    (3 inputs)
//  syndrom[38]:             x      x                         x   (3 inputs)
//  syndrom[39]:              x    x                         x    (3 inputs)
//  syndrom[40]:              x    x                          x   (3 inputs)
//  syndrom[41]:              x     x                        x    (3 inputs)
//  syndrom[42]:               x x                              x (3 inputs)
//  syndrom[43]:               x  x                            x  (3 inputs)
//  syndrom[44]:               x  x                             x (3 inputs)
//  syndrom[45]:                xx                             x  (3 inputs)
//  syndrom[46]:                xx                              x (3 inputs)
//  syndrom[47]:                x x                            x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 42 45 46)
//  input bit 17 used  3 times (syndrom bits 43 44 47)
//  input bit 18 used  3 times (syndrom bits 36 39 40)
//  input bit 19 used  3 times (syndrom bits 37 38 41)
//  input bit 20 used  3 times (syndrom bits 30 33 34)
//  input bit 21 used  3 times (syndrom bits 31 32 35)
//  input bit 22 used  3 times (syndrom bits 24 27 28)
//  input bit 23 used  3 times (syndrom bits 25 26 29)
//  input bit 24 used  3 times (syndrom bits 18 21 22)
//  input bit 25 used  3 times (syndrom bits 19 20 23)
//  input bit 26 used  3 times (syndrom bits 12 15 16)
//  input bit 27 used  3 times (syndrom bits 13 14 17)
//  input bit 28 used  3 times (syndrom bits 6 9 10)
//  input bit 29 used  3 times (syndrom bits 7 8 11)
//  input bit 30 used  3 times (syndrom bits 0 3 4)
//  input bit 31 used  3 times (syndrom bits 1 2 5)
//  input bit 32 used  3 times (syndrom bits 1 3 5)
//  input bit 33 used  3 times (syndrom bits 0 2 4)
//  input bit 34 used  3 times (syndrom bits 7 9 11)
//  input bit 35 used  3 times (syndrom bits 6 8 10)
//  input bit 36 used  3 times (syndrom bits 13 15 17)
//  input bit 37 used  3 times (syndrom bits 12 14 16)
//  input bit 38 used  3 times (syndrom bits 19 21 23)
//  input bit 39 used  3 times (syndrom bits 18 20 22)
//  input bit 40 used  3 times (syndrom bits 25 27 29)
//  input bit 41 used  3 times (syndrom bits 24 26 28)
//  input bit 42 used  3 times (syndrom bits 31 33 35)
//  input bit 43 used  3 times (syndrom bits 30 32 34)
//  input bit 44 used  3 times (syndrom bits 37 39 41)
//  input bit 45 used  3 times (syndrom bits 36 38 40)
//  input bit 46 used  3 times (syndrom bits 43 45 47)
//  input bit 47 used  3 times (syndrom bits 42 44 46)
function [48-1:0] extended_hamming_code_96_48_f;
    input [48-1:0] in;
    reg [48-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[30]^in[33];//3 inputs
        syndrom[ 1] = in[ 0]^in[31]^in[32];//3 inputs
        syndrom[ 2] = in[ 0]^in[31]^in[33];//3 inputs
        syndrom[ 3] = in[ 1]^in[30]^in[32];//3 inputs
        syndrom[ 4] = in[ 1]^in[30]^in[33];//3 inputs
        syndrom[ 5] = in[ 1]^in[31]^in[32];//3 inputs
        syndrom[ 6] = in[ 2]^in[28]^in[35];//3 inputs
        syndrom[ 7] = in[ 2]^in[29]^in[34];//3 inputs
        syndrom[ 8] = in[ 2]^in[29]^in[35];//3 inputs
        syndrom[ 9] = in[ 3]^in[28]^in[34];//3 inputs
        syndrom[10] = in[ 3]^in[28]^in[35];//3 inputs
        syndrom[11] = in[ 3]^in[29]^in[34];//3 inputs
        syndrom[12] = in[ 4]^in[26]^in[37];//3 inputs
        syndrom[13] = in[ 4]^in[27]^in[36];//3 inputs
        syndrom[14] = in[ 4]^in[27]^in[37];//3 inputs
        syndrom[15] = in[ 5]^in[26]^in[36];//3 inputs
        syndrom[16] = in[ 5]^in[26]^in[37];//3 inputs
        syndrom[17] = in[ 5]^in[27]^in[36];//3 inputs
        syndrom[18] = in[ 6]^in[24]^in[39];//3 inputs
        syndrom[19] = in[ 6]^in[25]^in[38];//3 inputs
        syndrom[20] = in[ 6]^in[25]^in[39];//3 inputs
        syndrom[21] = in[ 7]^in[24]^in[38];//3 inputs
        syndrom[22] = in[ 7]^in[24]^in[39];//3 inputs
        syndrom[23] = in[ 7]^in[25]^in[38];//3 inputs
        syndrom[24] = in[ 8]^in[22]^in[41];//3 inputs
        syndrom[25] = in[ 8]^in[23]^in[40];//3 inputs
        syndrom[26] = in[ 8]^in[23]^in[41];//3 inputs
        syndrom[27] = in[ 9]^in[22]^in[40];//3 inputs
        syndrom[28] = in[ 9]^in[22]^in[41];//3 inputs
        syndrom[29] = in[ 9]^in[23]^in[40];//3 inputs
        syndrom[30] = in[10]^in[20]^in[43];//3 inputs
        syndrom[31] = in[10]^in[21]^in[42];//3 inputs
        syndrom[32] = in[10]^in[21]^in[43];//3 inputs
        syndrom[33] = in[11]^in[20]^in[42];//3 inputs
        syndrom[34] = in[11]^in[20]^in[43];//3 inputs
        syndrom[35] = in[11]^in[21]^in[42];//3 inputs
        syndrom[36] = in[12]^in[18]^in[45];//3 inputs
        syndrom[37] = in[12]^in[19]^in[44];//3 inputs
        syndrom[38] = in[12]^in[19]^in[45];//3 inputs
        syndrom[39] = in[13]^in[18]^in[44];//3 inputs
        syndrom[40] = in[13]^in[18]^in[45];//3 inputs
        syndrom[41] = in[13]^in[19]^in[44];//3 inputs
        syndrom[42] = in[14]^in[16]^in[47];//3 inputs
        syndrom[43] = in[14]^in[17]^in[46];//3 inputs
        syndrom[44] = in[14]^in[17]^in[47];//3 inputs
        syndrom[45] = in[15]^in[16]^in[46];//3 inputs
        syndrom[46] = in[15]^in[16]^in[47];//3 inputs
        syndrom[47] = in[15]^in[17]^in[46];//3 inputs
        extended_hamming_code_96_48_f = syndrom;
    end
endfunction
function [2+48-1:0] extended_hamming_code_96_48_f_correction_pattern_f;
    input [48-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [48-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {48{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			48'b000000000000000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {48{1'b0}};
			end	
			48'b000000000000000000000000000000000000000000000111: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 0]=1'b1;
			end
			48'b000000000000000000000000000000000000000000111000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 1]=1'b1;
			end
			48'b000000000000000000000000000000000000000111000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 2]=1'b1;
			end
			48'b000000000000000000000000000000000000111000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 3]=1'b1;
			end
			48'b000000000000000000000000000000000111000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 4]=1'b1;
			end
			48'b000000000000000000000000000000111000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 5]=1'b1;
			end
			48'b000000000000000000000000000111000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 6]=1'b1;
			end
			48'b000000000000000000000000111000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 7]=1'b1;
			end
			48'b000000000000000000000111000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 8]=1'b1;
			end
			48'b000000000000000000111000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 9]=1'b1;
			end
			48'b000000000000000111000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[10]=1'b1;
			end
			48'b000000000000111000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[11]=1'b1;
			end
			48'b000000000111000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[12]=1'b1;
			end
			48'b000000111000000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[13]=1'b1;
			end
			48'b000111000000000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[14]=1'b1;
			end
			48'b111000000000000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[15]=1'b1;
			end
			48'b011001000000000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[16]=1'b1;
			end
			48'b100110000000000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[17]=1'b1;
			end
			48'b000000011001000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[18]=1'b1;
			end
			48'b000000100110000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[19]=1'b1;
			end
			48'b000000000000011001000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[20]=1'b1;
			end
			48'b000000000000100110000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[21]=1'b1;
			end
			48'b000000000000000000011001000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[22]=1'b1;
			end
			48'b000000000000000000100110000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[23]=1'b1;
			end
			48'b000000000000000000000000011001000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[24]=1'b1;
			end
			48'b000000000000000000000000100110000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[25]=1'b1;
			end
			48'b000000000000000000000000000000011001000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[26]=1'b1;
			end
			48'b000000000000000000000000000000100110000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[27]=1'b1;
			end
			48'b000000000000000000000000000000000000011001000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[28]=1'b1;
			end
			48'b000000000000000000000000000000000000100110000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[29]=1'b1;
			end
			48'b000000000000000000000000000000000000000000011001: begin
				correction_pattern = {48{1'b0}};correction_pattern[30]=1'b1;
			end
			48'b000000000000000000000000000000000000000000100110: begin
				correction_pattern = {48{1'b0}};correction_pattern[31]=1'b1;
			end
			48'b000000000000000000000000000000000000000000101010: begin
				correction_pattern = {48{1'b0}};correction_pattern[32]=1'b1;
			end
			48'b000000000000000000000000000000000000000000010101: begin
				correction_pattern = {48{1'b0}};correction_pattern[33]=1'b1;
			end
			48'b000000000000000000000000000000000000101010000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[34]=1'b1;
			end
			48'b000000000000000000000000000000000000010101000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[35]=1'b1;
			end
			48'b000000000000000000000000000000101010000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[36]=1'b1;
			end
			48'b000000000000000000000000000000010101000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[37]=1'b1;
			end
			48'b000000000000000000000000101010000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[38]=1'b1;
			end
			48'b000000000000000000000000010101000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[39]=1'b1;
			end
			48'b000000000000000000101010000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[40]=1'b1;
			end
			48'b000000000000000000010101000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[41]=1'b1;
			end
			48'b000000000000101010000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[42]=1'b1;
			end
			48'b000000000000010101000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[43]=1'b1;
			end
			48'b000000101010000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[44]=1'b1;
			end
			48'b000000010101000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[45]=1'b1;
			end
			48'b101010000000000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[46]=1'b1;
			end
			48'b010101000000000000000000000000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[47]=1'b1;
			end
			48'b000000000000000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000001000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000010000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000100000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000001000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000010000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000100000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000001000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000010000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000100000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b001000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b010000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b100000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_96_48_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [48-1:0] stored_data_edc = extended_hamming_code_96_48_f(i_stored_data);
wire [48-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [48-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_96_48_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_64_min_delay (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [64-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [64-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_128_64_f
//Compute 64 bits Error Detection Code from a 64 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 340282366920938463463374607431768211456 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[ 0]: x                                                             x  (2 inputs)
//  syndrom[ 1]: x                                                              x (2 inputs)
//  syndrom[ 2]:  x                                                            x  (2 inputs)
//  syndrom[ 3]:  x                                                             x (2 inputs)
//  syndrom[ 4]:   x                                                         x    (2 inputs)
//  syndrom[ 5]:   x                                                          x   (2 inputs)
//  syndrom[ 6]:    x                                                        x    (2 inputs)
//  syndrom[ 7]:    x                                                         x   (2 inputs)
//  syndrom[ 8]:     x                                                     x      (2 inputs)
//  syndrom[ 9]:     x                                                      x     (2 inputs)
//  syndrom[10]:      x                                                    x      (2 inputs)
//  syndrom[11]:      x                                                     x     (2 inputs)
//  syndrom[12]:       x                                                 x        (2 inputs)
//  syndrom[13]:       x                                                  x       (2 inputs)
//  syndrom[14]:        x                                                x        (2 inputs)
//  syndrom[15]:        x                                                 x       (2 inputs)
//  syndrom[16]:         x                                             x          (2 inputs)
//  syndrom[17]:         x                                              x         (2 inputs)
//  syndrom[18]:          x                                            x          (2 inputs)
//  syndrom[19]:          x                                             x         (2 inputs)
//  syndrom[20]:           x                                         x            (2 inputs)
//  syndrom[21]:           x                                          x           (2 inputs)
//  syndrom[22]:            x                                        x            (2 inputs)
//  syndrom[23]:            x                                         x           (2 inputs)
//  syndrom[24]:             x                                     x              (2 inputs)
//  syndrom[25]:             x                                      x             (2 inputs)
//  syndrom[26]:              x                                    x              (2 inputs)
//  syndrom[27]:              x                                     x             (2 inputs)
//  syndrom[28]:               x                                 x                (2 inputs)
//  syndrom[29]:               x                                  x               (2 inputs)
//  syndrom[30]:                x                                x                (2 inputs)
//  syndrom[31]:                x                                 x               (2 inputs)
//  syndrom[32]:                 x                             x                  (2 inputs)
//  syndrom[33]:                 x                              x                 (2 inputs)
//  syndrom[34]:                  x                            x                  (2 inputs)
//  syndrom[35]:                  x                             x                 (2 inputs)
//  syndrom[36]:                   x                         x                    (2 inputs)
//  syndrom[37]:                   x                          x                   (2 inputs)
//  syndrom[38]:                    x                        x                    (2 inputs)
//  syndrom[39]:                    x                         x                   (2 inputs)
//  syndrom[40]:                     x                     x                      (2 inputs)
//  syndrom[41]:                     x                      x                     (2 inputs)
//  syndrom[42]:                      x                    x                      (2 inputs)
//  syndrom[43]:                      x                     x                     (2 inputs)
//  syndrom[44]:                       x                 x                        (2 inputs)
//  syndrom[45]:                       x                  x                       (2 inputs)
//  syndrom[46]:                        x                x                        (2 inputs)
//  syndrom[47]:                        x                 x                       (2 inputs)
//  syndrom[48]:                         x             x                          (2 inputs)
//  syndrom[49]:                         x              x                         (2 inputs)
//  syndrom[50]:                          x            x                          (2 inputs)
//  syndrom[51]:                          x             x                         (2 inputs)
//  syndrom[52]:                           x         x                            (2 inputs)
//  syndrom[53]:                           x          x                           (2 inputs)
//  syndrom[54]:                            x        x                            (2 inputs)
//  syndrom[55]:                            x         x                           (2 inputs)
//  syndrom[56]:                             x     x                              (2 inputs)
//  syndrom[57]:                             x      x                             (2 inputs)
//  syndrom[58]:                              x    x                              (2 inputs)
//  syndrom[59]:                              x     x                             (2 inputs)
//  syndrom[60]:                               x x                                (2 inputs)
//  syndrom[61]:                               x  x                               (2 inputs)
//  syndrom[62]:                                xx                                (2 inputs)
//  syndrom[63]:                                x x                               (2 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 32 33)
//  input bit 17 used  2 times (syndrom bits 34 35)
//  input bit 18 used  2 times (syndrom bits 36 37)
//  input bit 19 used  2 times (syndrom bits 38 39)
//  input bit 20 used  2 times (syndrom bits 40 41)
//  input bit 21 used  2 times (syndrom bits 42 43)
//  input bit 22 used  2 times (syndrom bits 44 45)
//  input bit 23 used  2 times (syndrom bits 46 47)
//  input bit 24 used  2 times (syndrom bits 48 49)
//  input bit 25 used  2 times (syndrom bits 50 51)
//  input bit 26 used  2 times (syndrom bits 52 53)
//  input bit 27 used  2 times (syndrom bits 54 55)
//  input bit 28 used  2 times (syndrom bits 56 57)
//  input bit 29 used  2 times (syndrom bits 58 59)
//  input bit 30 used  2 times (syndrom bits 60 61)
//  input bit 31 used  2 times (syndrom bits 62 63)
//  input bit 32 used  2 times (syndrom bits 60 62)
//  input bit 33 used  2 times (syndrom bits 61 63)
//  input bit 34 used  2 times (syndrom bits 56 58)
//  input bit 35 used  2 times (syndrom bits 57 59)
//  input bit 36 used  2 times (syndrom bits 52 54)
//  input bit 37 used  2 times (syndrom bits 53 55)
//  input bit 38 used  2 times (syndrom bits 48 50)
//  input bit 39 used  2 times (syndrom bits 49 51)
//  input bit 40 used  2 times (syndrom bits 44 46)
//  input bit 41 used  2 times (syndrom bits 45 47)
//  input bit 42 used  2 times (syndrom bits 40 42)
//  input bit 43 used  2 times (syndrom bits 41 43)
//  input bit 44 used  2 times (syndrom bits 36 38)
//  input bit 45 used  2 times (syndrom bits 37 39)
//  input bit 46 used  2 times (syndrom bits 32 34)
//  input bit 47 used  2 times (syndrom bits 33 35)
//  input bit 48 used  2 times (syndrom bits 28 30)
//  input bit 49 used  2 times (syndrom bits 29 31)
//  input bit 50 used  2 times (syndrom bits 24 26)
//  input bit 51 used  2 times (syndrom bits 25 27)
//  input bit 52 used  2 times (syndrom bits 20 22)
//  input bit 53 used  2 times (syndrom bits 21 23)
//  input bit 54 used  2 times (syndrom bits 16 18)
//  input bit 55 used  2 times (syndrom bits 17 19)
//  input bit 56 used  2 times (syndrom bits 12 14)
//  input bit 57 used  2 times (syndrom bits 13 15)
//  input bit 58 used  2 times (syndrom bits 8 10)
//  input bit 59 used  2 times (syndrom bits 9 11)
//  input bit 60 used  2 times (syndrom bits 4 6)
//  input bit 61 used  2 times (syndrom bits 5 7)
//  input bit 62 used  2 times (syndrom bits 0 2)
//  input bit 63 used  2 times (syndrom bits 1 3)
function [64-1:0] hamming_code_128_64_f;
    input [64-1:0] in;
    reg [64-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[62];//2 inputs
        syndrom[ 1] = in[ 0]^in[63];//2 inputs
        syndrom[ 2] = in[ 1]^in[62];//2 inputs
        syndrom[ 3] = in[ 1]^in[63];//2 inputs
        syndrom[ 4] = in[ 2]^in[60];//2 inputs
        syndrom[ 5] = in[ 2]^in[61];//2 inputs
        syndrom[ 6] = in[ 3]^in[60];//2 inputs
        syndrom[ 7] = in[ 3]^in[61];//2 inputs
        syndrom[ 8] = in[ 4]^in[58];//2 inputs
        syndrom[ 9] = in[ 4]^in[59];//2 inputs
        syndrom[10] = in[ 5]^in[58];//2 inputs
        syndrom[11] = in[ 5]^in[59];//2 inputs
        syndrom[12] = in[ 6]^in[56];//2 inputs
        syndrom[13] = in[ 6]^in[57];//2 inputs
        syndrom[14] = in[ 7]^in[56];//2 inputs
        syndrom[15] = in[ 7]^in[57];//2 inputs
        syndrom[16] = in[ 8]^in[54];//2 inputs
        syndrom[17] = in[ 8]^in[55];//2 inputs
        syndrom[18] = in[ 9]^in[54];//2 inputs
        syndrom[19] = in[ 9]^in[55];//2 inputs
        syndrom[20] = in[10]^in[52];//2 inputs
        syndrom[21] = in[10]^in[53];//2 inputs
        syndrom[22] = in[11]^in[52];//2 inputs
        syndrom[23] = in[11]^in[53];//2 inputs
        syndrom[24] = in[12]^in[50];//2 inputs
        syndrom[25] = in[12]^in[51];//2 inputs
        syndrom[26] = in[13]^in[50];//2 inputs
        syndrom[27] = in[13]^in[51];//2 inputs
        syndrom[28] = in[14]^in[48];//2 inputs
        syndrom[29] = in[14]^in[49];//2 inputs
        syndrom[30] = in[15]^in[48];//2 inputs
        syndrom[31] = in[15]^in[49];//2 inputs
        syndrom[32] = in[16]^in[46];//2 inputs
        syndrom[33] = in[16]^in[47];//2 inputs
        syndrom[34] = in[17]^in[46];//2 inputs
        syndrom[35] = in[17]^in[47];//2 inputs
        syndrom[36] = in[18]^in[44];//2 inputs
        syndrom[37] = in[18]^in[45];//2 inputs
        syndrom[38] = in[19]^in[44];//2 inputs
        syndrom[39] = in[19]^in[45];//2 inputs
        syndrom[40] = in[20]^in[42];//2 inputs
        syndrom[41] = in[20]^in[43];//2 inputs
        syndrom[42] = in[21]^in[42];//2 inputs
        syndrom[43] = in[21]^in[43];//2 inputs
        syndrom[44] = in[22]^in[40];//2 inputs
        syndrom[45] = in[22]^in[41];//2 inputs
        syndrom[46] = in[23]^in[40];//2 inputs
        syndrom[47] = in[23]^in[41];//2 inputs
        syndrom[48] = in[24]^in[38];//2 inputs
        syndrom[49] = in[24]^in[39];//2 inputs
        syndrom[50] = in[25]^in[38];//2 inputs
        syndrom[51] = in[25]^in[39];//2 inputs
        syndrom[52] = in[26]^in[36];//2 inputs
        syndrom[53] = in[26]^in[37];//2 inputs
        syndrom[54] = in[27]^in[36];//2 inputs
        syndrom[55] = in[27]^in[37];//2 inputs
        syndrom[56] = in[28]^in[34];//2 inputs
        syndrom[57] = in[28]^in[35];//2 inputs
        syndrom[58] = in[29]^in[34];//2 inputs
        syndrom[59] = in[29]^in[35];//2 inputs
        syndrom[60] = in[30]^in[32];//2 inputs
        syndrom[61] = in[30]^in[33];//2 inputs
        syndrom[62] = in[31]^in[32];//2 inputs
        syndrom[63] = in[31]^in[33];//2 inputs
        hamming_code_128_64_f = syndrom;
    end
endfunction
wire [64-1:0] stored_data_edc = hamming_code_128_64_f(i_stored_data);
wire [64-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_64_min_delay (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [64-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [64-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_128_64_f
//Compute 64 bits Error Detection Code from a 64 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 340282366920938463463374607431768211456 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[ 0]: x                                        x  x                    (3 inputs)
//  syndrom[ 1]: x                                         xx                     (3 inputs)
//  syndrom[ 2]: x                                         xx                     (3 inputs)
//  syndrom[ 3]:  x                                      x    x                   (3 inputs)
//  syndrom[ 4]:  x                                       xx                      (3 inputs)
//  syndrom[ 5]:  x                                       x x                     (3 inputs)
//  syndrom[ 6]:   x                                    x      x                  (3 inputs)
//  syndrom[ 7]:   x                                     x   x                    (3 inputs)
//  syndrom[ 8]:   x                                     x   x                    (3 inputs)
//  syndrom[ 9]:    x                                  x        x                 (3 inputs)
//  syndrom[10]:    x                                   x     x                   (3 inputs)
//  syndrom[11]:    x                                   x     x                   (3 inputs)
//  syndrom[12]:     x                                x          x                (3 inputs)
//  syndrom[13]:     x                                 x       x                  (3 inputs)
//  syndrom[14]:     x                                 x       x                  (3 inputs)
//  syndrom[15]:      x                              x            x               (3 inputs)
//  syndrom[16]:      x                               x         x                 (3 inputs)
//  syndrom[17]:      x                               x         x                 (3 inputs)
//  syndrom[18]:       x                            x              x              (3 inputs)
//  syndrom[19]:       x                             x           x                (3 inputs)
//  syndrom[20]:       x                             x           x                (3 inputs)
//  syndrom[21]:        x                          x                x             (3 inputs)
//  syndrom[22]:        x                           x             x               (3 inputs)
//  syndrom[23]:        x                           x             x               (3 inputs)
//  syndrom[24]:         x                        x                  x            (3 inputs)
//  syndrom[25]:         x                         x               x              (3 inputs)
//  syndrom[26]:         x                         x               x              (3 inputs)
//  syndrom[27]:          x                      x                    x           (3 inputs)
//  syndrom[28]:          x                       x                 x             (3 inputs)
//  syndrom[29]:          x                       x                 x             (3 inputs)
//  syndrom[30]:           x                    x                      x          (3 inputs)
//  syndrom[31]:           x                     x                   x            (3 inputs)
//  syndrom[32]:           x                     x                   x            (3 inputs)
//  syndrom[33]:            x                  x                        x         (3 inputs)
//  syndrom[34]:            x                   x                     x           (3 inputs)
//  syndrom[35]:            x                   x                     x           (3 inputs)
//  syndrom[36]:             x                x                          x        (3 inputs)
//  syndrom[37]:             x                 x                       x          (3 inputs)
//  syndrom[38]:             x                 x                       x          (3 inputs)
//  syndrom[39]:              x              x                            x       (3 inputs)
//  syndrom[40]:              x               x                         x         (3 inputs)
//  syndrom[41]:              x               x                         x         (3 inputs)
//  syndrom[42]:               x            x                              x      (3 inputs)
//  syndrom[43]:               x             x                           x        (3 inputs)
//  syndrom[44]:               x             x                           x        (3 inputs)
//  syndrom[45]:                x          x                                x     (3 inputs)
//  syndrom[46]:                x           x                             x       (3 inputs)
//  syndrom[47]:                x           x                             x       (3 inputs)
//  syndrom[48]:                 x        x                                  x    (3 inputs)
//  syndrom[49]:                 x         x                               x      (3 inputs)
//  syndrom[50]:                 x         x                               x      (3 inputs)
//  syndrom[51]:                  x      x                                    x   (3 inputs)
//  syndrom[52]:                  x       x                                 x     (3 inputs)
//  syndrom[53]:                  x       x                                 x     (3 inputs)
//  syndrom[54]:                   x    x                                      x  (3 inputs)
//  syndrom[55]:                   x     x                                   x    (3 inputs)
//  syndrom[56]:                   x     x                                   x    (3 inputs)
//  syndrom[57]:                    x  x                                        x (3 inputs)
//  syndrom[58]:                    x   x                                     x   (3 inputs)
//  syndrom[59]:                    x   x                                     x   (3 inputs)
//  syndrom[60]:                     xx                                         x (3 inputs)
//  syndrom[61]:                     xx                                         x (3 inputs)
//  syndrom[62]:                     x x                                       x  (3 inputs)
//  syndrom[63]:                      xx                                       x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 48 49 50)
//  input bit 17 used  3 times (syndrom bits 51 52 53)
//  input bit 18 used  3 times (syndrom bits 54 55 56)
//  input bit 19 used  3 times (syndrom bits 57 58 59)
//  input bit 20 used  3 times (syndrom bits 60 61 62)
//  input bit 21 used  3 times (syndrom bits 60 61 63)
//  input bit 22 used  3 times (syndrom bits 57 62 63)
//  input bit 23 used  3 times (syndrom bits 54 58 59)
//  input bit 24 used  3 times (syndrom bits 51 55 56)
//  input bit 25 used  3 times (syndrom bits 48 52 53)
//  input bit 26 used  3 times (syndrom bits 45 49 50)
//  input bit 27 used  3 times (syndrom bits 42 46 47)
//  input bit 28 used  3 times (syndrom bits 39 43 44)
//  input bit 29 used  3 times (syndrom bits 36 40 41)
//  input bit 30 used  3 times (syndrom bits 33 37 38)
//  input bit 31 used  3 times (syndrom bits 30 34 35)
//  input bit 32 used  3 times (syndrom bits 27 31 32)
//  input bit 33 used  3 times (syndrom bits 24 28 29)
//  input bit 34 used  3 times (syndrom bits 21 25 26)
//  input bit 35 used  3 times (syndrom bits 18 22 23)
//  input bit 36 used  3 times (syndrom bits 15 19 20)
//  input bit 37 used  3 times (syndrom bits 12 16 17)
//  input bit 38 used  3 times (syndrom bits 9 13 14)
//  input bit 39 used  3 times (syndrom bits 6 10 11)
//  input bit 40 used  3 times (syndrom bits 3 7 8)
//  input bit 41 used  3 times (syndrom bits 0 4 5)
//  input bit 42 used  3 times (syndrom bits 1 2 4)
//  input bit 43 used  3 times (syndrom bits 1 2 5)
//  input bit 44 used  3 times (syndrom bits 0 7 8)
//  input bit 45 used  3 times (syndrom bits 3 10 11)
//  input bit 46 used  3 times (syndrom bits 6 13 14)
//  input bit 47 used  3 times (syndrom bits 9 16 17)
//  input bit 48 used  3 times (syndrom bits 12 19 20)
//  input bit 49 used  3 times (syndrom bits 15 22 23)
//  input bit 50 used  3 times (syndrom bits 18 25 26)
//  input bit 51 used  3 times (syndrom bits 21 28 29)
//  input bit 52 used  3 times (syndrom bits 24 31 32)
//  input bit 53 used  3 times (syndrom bits 27 34 35)
//  input bit 54 used  3 times (syndrom bits 30 37 38)
//  input bit 55 used  3 times (syndrom bits 33 40 41)
//  input bit 56 used  3 times (syndrom bits 36 43 44)
//  input bit 57 used  3 times (syndrom bits 39 46 47)
//  input bit 58 used  3 times (syndrom bits 42 49 50)
//  input bit 59 used  3 times (syndrom bits 45 52 53)
//  input bit 60 used  3 times (syndrom bits 48 55 56)
//  input bit 61 used  3 times (syndrom bits 51 58 59)
//  input bit 62 used  3 times (syndrom bits 54 62 63)
//  input bit 63 used  3 times (syndrom bits 57 60 61)
function [64-1:0] extended_hamming_code_128_64_f;
    input [64-1:0] in;
    reg [64-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[41]^in[44];//3 inputs
        syndrom[ 1] = in[ 0]^in[42]^in[43];//3 inputs
        syndrom[ 2] = in[ 0]^in[42]^in[43];//3 inputs
        syndrom[ 3] = in[ 1]^in[40]^in[45];//3 inputs
        syndrom[ 4] = in[ 1]^in[41]^in[42];//3 inputs
        syndrom[ 5] = in[ 1]^in[41]^in[43];//3 inputs
        syndrom[ 6] = in[ 2]^in[39]^in[46];//3 inputs
        syndrom[ 7] = in[ 2]^in[40]^in[44];//3 inputs
        syndrom[ 8] = in[ 2]^in[40]^in[44];//3 inputs
        syndrom[ 9] = in[ 3]^in[38]^in[47];//3 inputs
        syndrom[10] = in[ 3]^in[39]^in[45];//3 inputs
        syndrom[11] = in[ 3]^in[39]^in[45];//3 inputs
        syndrom[12] = in[ 4]^in[37]^in[48];//3 inputs
        syndrom[13] = in[ 4]^in[38]^in[46];//3 inputs
        syndrom[14] = in[ 4]^in[38]^in[46];//3 inputs
        syndrom[15] = in[ 5]^in[36]^in[49];//3 inputs
        syndrom[16] = in[ 5]^in[37]^in[47];//3 inputs
        syndrom[17] = in[ 5]^in[37]^in[47];//3 inputs
        syndrom[18] = in[ 6]^in[35]^in[50];//3 inputs
        syndrom[19] = in[ 6]^in[36]^in[48];//3 inputs
        syndrom[20] = in[ 6]^in[36]^in[48];//3 inputs
        syndrom[21] = in[ 7]^in[34]^in[51];//3 inputs
        syndrom[22] = in[ 7]^in[35]^in[49];//3 inputs
        syndrom[23] = in[ 7]^in[35]^in[49];//3 inputs
        syndrom[24] = in[ 8]^in[33]^in[52];//3 inputs
        syndrom[25] = in[ 8]^in[34]^in[50];//3 inputs
        syndrom[26] = in[ 8]^in[34]^in[50];//3 inputs
        syndrom[27] = in[ 9]^in[32]^in[53];//3 inputs
        syndrom[28] = in[ 9]^in[33]^in[51];//3 inputs
        syndrom[29] = in[ 9]^in[33]^in[51];//3 inputs
        syndrom[30] = in[10]^in[31]^in[54];//3 inputs
        syndrom[31] = in[10]^in[32]^in[52];//3 inputs
        syndrom[32] = in[10]^in[32]^in[52];//3 inputs
        syndrom[33] = in[11]^in[30]^in[55];//3 inputs
        syndrom[34] = in[11]^in[31]^in[53];//3 inputs
        syndrom[35] = in[11]^in[31]^in[53];//3 inputs
        syndrom[36] = in[12]^in[29]^in[56];//3 inputs
        syndrom[37] = in[12]^in[30]^in[54];//3 inputs
        syndrom[38] = in[12]^in[30]^in[54];//3 inputs
        syndrom[39] = in[13]^in[28]^in[57];//3 inputs
        syndrom[40] = in[13]^in[29]^in[55];//3 inputs
        syndrom[41] = in[13]^in[29]^in[55];//3 inputs
        syndrom[42] = in[14]^in[27]^in[58];//3 inputs
        syndrom[43] = in[14]^in[28]^in[56];//3 inputs
        syndrom[44] = in[14]^in[28]^in[56];//3 inputs
        syndrom[45] = in[15]^in[26]^in[59];//3 inputs
        syndrom[46] = in[15]^in[27]^in[57];//3 inputs
        syndrom[47] = in[15]^in[27]^in[57];//3 inputs
        syndrom[48] = in[16]^in[25]^in[60];//3 inputs
        syndrom[49] = in[16]^in[26]^in[58];//3 inputs
        syndrom[50] = in[16]^in[26]^in[58];//3 inputs
        syndrom[51] = in[17]^in[24]^in[61];//3 inputs
        syndrom[52] = in[17]^in[25]^in[59];//3 inputs
        syndrom[53] = in[17]^in[25]^in[59];//3 inputs
        syndrom[54] = in[18]^in[23]^in[62];//3 inputs
        syndrom[55] = in[18]^in[24]^in[60];//3 inputs
        syndrom[56] = in[18]^in[24]^in[60];//3 inputs
        syndrom[57] = in[19]^in[22]^in[63];//3 inputs
        syndrom[58] = in[19]^in[23]^in[61];//3 inputs
        syndrom[59] = in[19]^in[23]^in[61];//3 inputs
        syndrom[60] = in[20]^in[21]^in[63];//3 inputs
        syndrom[61] = in[20]^in[21]^in[63];//3 inputs
        syndrom[62] = in[20]^in[22]^in[62];//3 inputs
        syndrom[63] = in[21]^in[22]^in[62];//3 inputs
        extended_hamming_code_128_64_f = syndrom;
    end
endfunction
wire [64-1:0] stored_data_edc = extended_hamming_code_128_64_f(i_stored_data);
wire [64-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_64_min_delay (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [64-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [64-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [64-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_128_64_f
//Compute 64 bits Error Detection Code from a 64 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 340282366920938463463374607431768211456 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[ 0]: x                                        x  x                    (3 inputs)
//  syndrom[ 1]: x                                         xx                     (3 inputs)
//  syndrom[ 2]: x                                         xx                     (3 inputs)
//  syndrom[ 3]:  x                                      x    x                   (3 inputs)
//  syndrom[ 4]:  x                                       xx                      (3 inputs)
//  syndrom[ 5]:  x                                       x x                     (3 inputs)
//  syndrom[ 6]:   x                                    x      x                  (3 inputs)
//  syndrom[ 7]:   x                                     x   x                    (3 inputs)
//  syndrom[ 8]:   x                                     x   x                    (3 inputs)
//  syndrom[ 9]:    x                                  x        x                 (3 inputs)
//  syndrom[10]:    x                                   x     x                   (3 inputs)
//  syndrom[11]:    x                                   x     x                   (3 inputs)
//  syndrom[12]:     x                                x          x                (3 inputs)
//  syndrom[13]:     x                                 x       x                  (3 inputs)
//  syndrom[14]:     x                                 x       x                  (3 inputs)
//  syndrom[15]:      x                              x            x               (3 inputs)
//  syndrom[16]:      x                               x         x                 (3 inputs)
//  syndrom[17]:      x                               x         x                 (3 inputs)
//  syndrom[18]:       x                            x              x              (3 inputs)
//  syndrom[19]:       x                             x           x                (3 inputs)
//  syndrom[20]:       x                             x           x                (3 inputs)
//  syndrom[21]:        x                          x                x             (3 inputs)
//  syndrom[22]:        x                           x             x               (3 inputs)
//  syndrom[23]:        x                           x             x               (3 inputs)
//  syndrom[24]:         x                        x                  x            (3 inputs)
//  syndrom[25]:         x                         x               x              (3 inputs)
//  syndrom[26]:         x                         x               x              (3 inputs)
//  syndrom[27]:          x                      x                    x           (3 inputs)
//  syndrom[28]:          x                       x                 x             (3 inputs)
//  syndrom[29]:          x                       x                 x             (3 inputs)
//  syndrom[30]:           x                    x                      x          (3 inputs)
//  syndrom[31]:           x                     x                   x            (3 inputs)
//  syndrom[32]:           x                     x                   x            (3 inputs)
//  syndrom[33]:            x                  x                        x         (3 inputs)
//  syndrom[34]:            x                   x                     x           (3 inputs)
//  syndrom[35]:            x                   x                     x           (3 inputs)
//  syndrom[36]:             x                x                          x        (3 inputs)
//  syndrom[37]:             x                 x                       x          (3 inputs)
//  syndrom[38]:             x                 x                       x          (3 inputs)
//  syndrom[39]:              x              x                            x       (3 inputs)
//  syndrom[40]:              x               x                         x         (3 inputs)
//  syndrom[41]:              x               x                         x         (3 inputs)
//  syndrom[42]:               x            x                              x      (3 inputs)
//  syndrom[43]:               x             x                           x        (3 inputs)
//  syndrom[44]:               x             x                           x        (3 inputs)
//  syndrom[45]:                x          x                                x     (3 inputs)
//  syndrom[46]:                x           x                             x       (3 inputs)
//  syndrom[47]:                x           x                             x       (3 inputs)
//  syndrom[48]:                 x        x                                  x    (3 inputs)
//  syndrom[49]:                 x         x                               x      (3 inputs)
//  syndrom[50]:                 x         x                               x      (3 inputs)
//  syndrom[51]:                  x      x                                    x   (3 inputs)
//  syndrom[52]:                  x       x                                 x     (3 inputs)
//  syndrom[53]:                  x       x                                 x     (3 inputs)
//  syndrom[54]:                   x    x                                      x  (3 inputs)
//  syndrom[55]:                   x     x                                   x    (3 inputs)
//  syndrom[56]:                   x     x                                   x    (3 inputs)
//  syndrom[57]:                    x  x                                        x (3 inputs)
//  syndrom[58]:                    x   x                                     x   (3 inputs)
//  syndrom[59]:                    x   x                                     x   (3 inputs)
//  syndrom[60]:                     xx                                         x (3 inputs)
//  syndrom[61]:                     xx                                         x (3 inputs)
//  syndrom[62]:                     x x                                       x  (3 inputs)
//  syndrom[63]:                      xx                                       x  (3 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 48 49 50)
//  input bit 17 used  3 times (syndrom bits 51 52 53)
//  input bit 18 used  3 times (syndrom bits 54 55 56)
//  input bit 19 used  3 times (syndrom bits 57 58 59)
//  input bit 20 used  3 times (syndrom bits 60 61 62)
//  input bit 21 used  3 times (syndrom bits 60 61 63)
//  input bit 22 used  3 times (syndrom bits 57 62 63)
//  input bit 23 used  3 times (syndrom bits 54 58 59)
//  input bit 24 used  3 times (syndrom bits 51 55 56)
//  input bit 25 used  3 times (syndrom bits 48 52 53)
//  input bit 26 used  3 times (syndrom bits 45 49 50)
//  input bit 27 used  3 times (syndrom bits 42 46 47)
//  input bit 28 used  3 times (syndrom bits 39 43 44)
//  input bit 29 used  3 times (syndrom bits 36 40 41)
//  input bit 30 used  3 times (syndrom bits 33 37 38)
//  input bit 31 used  3 times (syndrom bits 30 34 35)
//  input bit 32 used  3 times (syndrom bits 27 31 32)
//  input bit 33 used  3 times (syndrom bits 24 28 29)
//  input bit 34 used  3 times (syndrom bits 21 25 26)
//  input bit 35 used  3 times (syndrom bits 18 22 23)
//  input bit 36 used  3 times (syndrom bits 15 19 20)
//  input bit 37 used  3 times (syndrom bits 12 16 17)
//  input bit 38 used  3 times (syndrom bits 9 13 14)
//  input bit 39 used  3 times (syndrom bits 6 10 11)
//  input bit 40 used  3 times (syndrom bits 3 7 8)
//  input bit 41 used  3 times (syndrom bits 0 4 5)
//  input bit 42 used  3 times (syndrom bits 1 2 4)
//  input bit 43 used  3 times (syndrom bits 1 2 5)
//  input bit 44 used  3 times (syndrom bits 0 7 8)
//  input bit 45 used  3 times (syndrom bits 3 10 11)
//  input bit 46 used  3 times (syndrom bits 6 13 14)
//  input bit 47 used  3 times (syndrom bits 9 16 17)
//  input bit 48 used  3 times (syndrom bits 12 19 20)
//  input bit 49 used  3 times (syndrom bits 15 22 23)
//  input bit 50 used  3 times (syndrom bits 18 25 26)
//  input bit 51 used  3 times (syndrom bits 21 28 29)
//  input bit 52 used  3 times (syndrom bits 24 31 32)
//  input bit 53 used  3 times (syndrom bits 27 34 35)
//  input bit 54 used  3 times (syndrom bits 30 37 38)
//  input bit 55 used  3 times (syndrom bits 33 40 41)
//  input bit 56 used  3 times (syndrom bits 36 43 44)
//  input bit 57 used  3 times (syndrom bits 39 46 47)
//  input bit 58 used  3 times (syndrom bits 42 49 50)
//  input bit 59 used  3 times (syndrom bits 45 52 53)
//  input bit 60 used  3 times (syndrom bits 48 55 56)
//  input bit 61 used  3 times (syndrom bits 51 58 59)
//  input bit 62 used  3 times (syndrom bits 54 62 63)
//  input bit 63 used  3 times (syndrom bits 57 60 61)
function [64-1:0] extended_hamming_code_128_64_f;
    input [64-1:0] in;
    reg [64-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[41]^in[44];//3 inputs
        syndrom[ 1] = in[ 0]^in[42]^in[43];//3 inputs
        syndrom[ 2] = in[ 0]^in[42]^in[43];//3 inputs
        syndrom[ 3] = in[ 1]^in[40]^in[45];//3 inputs
        syndrom[ 4] = in[ 1]^in[41]^in[42];//3 inputs
        syndrom[ 5] = in[ 1]^in[41]^in[43];//3 inputs
        syndrom[ 6] = in[ 2]^in[39]^in[46];//3 inputs
        syndrom[ 7] = in[ 2]^in[40]^in[44];//3 inputs
        syndrom[ 8] = in[ 2]^in[40]^in[44];//3 inputs
        syndrom[ 9] = in[ 3]^in[38]^in[47];//3 inputs
        syndrom[10] = in[ 3]^in[39]^in[45];//3 inputs
        syndrom[11] = in[ 3]^in[39]^in[45];//3 inputs
        syndrom[12] = in[ 4]^in[37]^in[48];//3 inputs
        syndrom[13] = in[ 4]^in[38]^in[46];//3 inputs
        syndrom[14] = in[ 4]^in[38]^in[46];//3 inputs
        syndrom[15] = in[ 5]^in[36]^in[49];//3 inputs
        syndrom[16] = in[ 5]^in[37]^in[47];//3 inputs
        syndrom[17] = in[ 5]^in[37]^in[47];//3 inputs
        syndrom[18] = in[ 6]^in[35]^in[50];//3 inputs
        syndrom[19] = in[ 6]^in[36]^in[48];//3 inputs
        syndrom[20] = in[ 6]^in[36]^in[48];//3 inputs
        syndrom[21] = in[ 7]^in[34]^in[51];//3 inputs
        syndrom[22] = in[ 7]^in[35]^in[49];//3 inputs
        syndrom[23] = in[ 7]^in[35]^in[49];//3 inputs
        syndrom[24] = in[ 8]^in[33]^in[52];//3 inputs
        syndrom[25] = in[ 8]^in[34]^in[50];//3 inputs
        syndrom[26] = in[ 8]^in[34]^in[50];//3 inputs
        syndrom[27] = in[ 9]^in[32]^in[53];//3 inputs
        syndrom[28] = in[ 9]^in[33]^in[51];//3 inputs
        syndrom[29] = in[ 9]^in[33]^in[51];//3 inputs
        syndrom[30] = in[10]^in[31]^in[54];//3 inputs
        syndrom[31] = in[10]^in[32]^in[52];//3 inputs
        syndrom[32] = in[10]^in[32]^in[52];//3 inputs
        syndrom[33] = in[11]^in[30]^in[55];//3 inputs
        syndrom[34] = in[11]^in[31]^in[53];//3 inputs
        syndrom[35] = in[11]^in[31]^in[53];//3 inputs
        syndrom[36] = in[12]^in[29]^in[56];//3 inputs
        syndrom[37] = in[12]^in[30]^in[54];//3 inputs
        syndrom[38] = in[12]^in[30]^in[54];//3 inputs
        syndrom[39] = in[13]^in[28]^in[57];//3 inputs
        syndrom[40] = in[13]^in[29]^in[55];//3 inputs
        syndrom[41] = in[13]^in[29]^in[55];//3 inputs
        syndrom[42] = in[14]^in[27]^in[58];//3 inputs
        syndrom[43] = in[14]^in[28]^in[56];//3 inputs
        syndrom[44] = in[14]^in[28]^in[56];//3 inputs
        syndrom[45] = in[15]^in[26]^in[59];//3 inputs
        syndrom[46] = in[15]^in[27]^in[57];//3 inputs
        syndrom[47] = in[15]^in[27]^in[57];//3 inputs
        syndrom[48] = in[16]^in[25]^in[60];//3 inputs
        syndrom[49] = in[16]^in[26]^in[58];//3 inputs
        syndrom[50] = in[16]^in[26]^in[58];//3 inputs
        syndrom[51] = in[17]^in[24]^in[61];//3 inputs
        syndrom[52] = in[17]^in[25]^in[59];//3 inputs
        syndrom[53] = in[17]^in[25]^in[59];//3 inputs
        syndrom[54] = in[18]^in[23]^in[62];//3 inputs
        syndrom[55] = in[18]^in[24]^in[60];//3 inputs
        syndrom[56] = in[18]^in[24]^in[60];//3 inputs
        syndrom[57] = in[19]^in[22]^in[63];//3 inputs
        syndrom[58] = in[19]^in[23]^in[61];//3 inputs
        syndrom[59] = in[19]^in[23]^in[61];//3 inputs
        syndrom[60] = in[20]^in[21]^in[63];//3 inputs
        syndrom[61] = in[20]^in[21]^in[63];//3 inputs
        syndrom[62] = in[20]^in[22]^in[62];//3 inputs
        syndrom[63] = in[21]^in[22]^in[62];//3 inputs
        extended_hamming_code_128_64_f = syndrom;
    end
endfunction
function [2+64-1:0] extended_hamming_code_128_64_f_correction_pattern_f;
    input [64-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [64-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {64{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			64'b0000000000000000000000000000000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {64{1'b0}};
			end	
			64'b0000000000000000000000000000000000000000000000000000000000000111: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 0]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000111000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 1]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000111000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 2]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000111000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 3]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000111000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 4]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000111000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 5]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000111000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 6]=1'b1;
			end
			64'b0000000000000000000000000000000000000000111000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 7]=1'b1;
			end
			64'b0000000000000000000000000000000000000111000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 8]=1'b1;
			end
			64'b0000000000000000000000000000000000111000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 9]=1'b1;
			end
			64'b0000000000000000000000000000000111000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[10]=1'b1;
			end
			64'b0000000000000000000000000000111000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[11]=1'b1;
			end
			64'b0000000000000000000000000111000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[12]=1'b1;
			end
			64'b0000000000000000000000111000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[13]=1'b1;
			end
			64'b0000000000000000000111000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[14]=1'b1;
			end
			64'b0000000000000000111000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[15]=1'b1;
			end
			64'b0000000000000111000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[16]=1'b1;
			end
			64'b0000000000111000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[17]=1'b1;
			end
			64'b0000000111000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[18]=1'b1;
			end
			64'b0000111000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[19]=1'b1;
			end
			64'b0111000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[20]=1'b1;
			end
			64'b1011000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[21]=1'b1;
			end
			64'b1100001000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[22]=1'b1;
			end
			64'b0000110001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[23]=1'b1;
			end
			64'b0000000110001000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[24]=1'b1;
			end
			64'b0000000000110001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[25]=1'b1;
			end
			64'b0000000000000110001000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[26]=1'b1;
			end
			64'b0000000000000000110001000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[27]=1'b1;
			end
			64'b0000000000000000000110001000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[28]=1'b1;
			end
			64'b0000000000000000000000110001000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[29]=1'b1;
			end
			64'b0000000000000000000000000110001000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[30]=1'b1;
			end
			64'b0000000000000000000000000000110001000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[31]=1'b1;
			end
			64'b0000000000000000000000000000000110001000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[32]=1'b1;
			end
			64'b0000000000000000000000000000000000110001000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[33]=1'b1;
			end
			64'b0000000000000000000000000000000000000110001000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[34]=1'b1;
			end
			64'b0000000000000000000000000000000000000000110001000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[35]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000110001000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[36]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000110001000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[37]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000110001000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[38]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000110001000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[39]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000110001000: begin
				correction_pattern = {64{1'b0}};correction_pattern[40]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000110001: begin
				correction_pattern = {64{1'b0}};correction_pattern[41]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000010110: begin
				correction_pattern = {64{1'b0}};correction_pattern[42]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000100110: begin
				correction_pattern = {64{1'b0}};correction_pattern[43]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000110000001: begin
				correction_pattern = {64{1'b0}};correction_pattern[44]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000110000001000: begin
				correction_pattern = {64{1'b0}};correction_pattern[45]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000110000001000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[46]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000110000001000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[47]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000110000001000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[48]=1'b1;
			end
			64'b0000000000000000000000000000000000000000110000001000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[49]=1'b1;
			end
			64'b0000000000000000000000000000000000000110000001000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[50]=1'b1;
			end
			64'b0000000000000000000000000000000000110000001000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[51]=1'b1;
			end
			64'b0000000000000000000000000000000110000001000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[52]=1'b1;
			end
			64'b0000000000000000000000000000110000001000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[53]=1'b1;
			end
			64'b0000000000000000000000000110000001000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[54]=1'b1;
			end
			64'b0000000000000000000000110000001000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[55]=1'b1;
			end
			64'b0000000000000000000110000001000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[56]=1'b1;
			end
			64'b0000000000000000110000001000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[57]=1'b1;
			end
			64'b0000000000000110000001000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[58]=1'b1;
			end
			64'b0000000000110000001000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[59]=1'b1;
			end
			64'b0000000110000001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[60]=1'b1;
			end
			64'b0000110000001000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[61]=1'b1;
			end
			64'b1100000001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[62]=1'b1;
			end
			64'b0011001000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[63]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000001000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000010000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000100000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000001000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000010000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000100000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000001000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000010000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000100000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000001000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000010000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000100000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000001000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000010000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000100000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000001000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000010000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000100000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000001000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000010000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000100000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000001000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000010000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000100000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0001000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0010000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0100000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b1000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_128_64_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [64-1:0] stored_data_edc = extended_hamming_code_128_64_f(i_stored_data);
wire [64-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [64-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_128_64_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_96_min_delay (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [96-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [96-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_192_96_f
//Compute 96 bits Error Detection Code from a 96 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 32 33)
//  input bit 17 used  2 times (syndrom bits 34 35)
//  input bit 18 used  2 times (syndrom bits 36 37)
//  input bit 19 used  2 times (syndrom bits 38 39)
//  input bit 20 used  2 times (syndrom bits 40 41)
//  input bit 21 used  2 times (syndrom bits 42 43)
//  input bit 22 used  2 times (syndrom bits 44 45)
//  input bit 23 used  2 times (syndrom bits 46 47)
//  input bit 24 used  2 times (syndrom bits 48 49)
//  input bit 25 used  2 times (syndrom bits 50 51)
//  input bit 26 used  2 times (syndrom bits 52 53)
//  input bit 27 used  2 times (syndrom bits 54 55)
//  input bit 28 used  2 times (syndrom bits 56 57)
//  input bit 29 used  2 times (syndrom bits 58 59)
//  input bit 30 used  2 times (syndrom bits 60 61)
//  input bit 31 used  2 times (syndrom bits 62 63)
//  input bit 32 used  2 times (syndrom bits 64 65)
//  input bit 33 used  2 times (syndrom bits 66 67)
//  input bit 34 used  2 times (syndrom bits 68 69)
//  input bit 35 used  2 times (syndrom bits 70 71)
//  input bit 36 used  2 times (syndrom bits 72 73)
//  input bit 37 used  2 times (syndrom bits 74 75)
//  input bit 38 used  2 times (syndrom bits 76 77)
//  input bit 39 used  2 times (syndrom bits 78 79)
//  input bit 40 used  2 times (syndrom bits 80 81)
//  input bit 41 used  2 times (syndrom bits 82 83)
//  input bit 42 used  2 times (syndrom bits 84 85)
//  input bit 43 used  2 times (syndrom bits 86 87)
//  input bit 44 used  2 times (syndrom bits 88 89)
//  input bit 45 used  2 times (syndrom bits 90 91)
//  input bit 46 used  2 times (syndrom bits 92 93)
//  input bit 47 used  2 times (syndrom bits 94 95)
//  input bit 48 used  2 times (syndrom bits 92 94)
//  input bit 49 used  2 times (syndrom bits 93 95)
//  input bit 50 used  2 times (syndrom bits 88 90)
//  input bit 51 used  2 times (syndrom bits 89 91)
//  input bit 52 used  2 times (syndrom bits 84 86)
//  input bit 53 used  2 times (syndrom bits 85 87)
//  input bit 54 used  2 times (syndrom bits 80 82)
//  input bit 55 used  2 times (syndrom bits 81 83)
//  input bit 56 used  2 times (syndrom bits 76 78)
//  input bit 57 used  2 times (syndrom bits 77 79)
//  input bit 58 used  2 times (syndrom bits 72 74)
//  input bit 59 used  2 times (syndrom bits 73 75)
//  input bit 60 used  2 times (syndrom bits 68 70)
//  input bit 61 used  2 times (syndrom bits 69 71)
//  input bit 62 used  2 times (syndrom bits 64 66)
//  input bit 63 used  2 times (syndrom bits 65 67)
//  input bit 64 used  2 times (syndrom bits 60 62)
//  input bit 65 used  2 times (syndrom bits 61 63)
//  input bit 66 used  2 times (syndrom bits 56 58)
//  input bit 67 used  2 times (syndrom bits 57 59)
//  input bit 68 used  2 times (syndrom bits 52 54)
//  input bit 69 used  2 times (syndrom bits 53 55)
//  input bit 70 used  2 times (syndrom bits 48 50)
//  input bit 71 used  2 times (syndrom bits 49 51)
//  input bit 72 used  2 times (syndrom bits 44 46)
//  input bit 73 used  2 times (syndrom bits 45 47)
//  input bit 74 used  2 times (syndrom bits 40 42)
//  input bit 75 used  2 times (syndrom bits 41 43)
//  input bit 76 used  2 times (syndrom bits 36 38)
//  input bit 77 used  2 times (syndrom bits 37 39)
//  input bit 78 used  2 times (syndrom bits 32 34)
//  input bit 79 used  2 times (syndrom bits 33 35)
//  input bit 80 used  2 times (syndrom bits 28 30)
//  input bit 81 used  2 times (syndrom bits 29 31)
//  input bit 82 used  2 times (syndrom bits 24 26)
//  input bit 83 used  2 times (syndrom bits 25 27)
//  input bit 84 used  2 times (syndrom bits 20 22)
//  input bit 85 used  2 times (syndrom bits 21 23)
//  input bit 86 used  2 times (syndrom bits 16 18)
//  input bit 87 used  2 times (syndrom bits 17 19)
//  input bit 88 used  2 times (syndrom bits 12 14)
//  input bit 89 used  2 times (syndrom bits 13 15)
//  input bit 90 used  2 times (syndrom bits 8 10)
//  input bit 91 used  2 times (syndrom bits 9 11)
//  input bit 92 used  2 times (syndrom bits 4 6)
//  input bit 93 used  2 times (syndrom bits 5 7)
//  input bit 94 used  2 times (syndrom bits 0 2)
//  input bit 95 used  2 times (syndrom bits 1 3)
function [96-1:0] hamming_code_192_96_f;
    input [96-1:0] in;
    reg [96-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[94];//2 inputs
        syndrom[ 1] = in[ 0]^in[95];//2 inputs
        syndrom[ 2] = in[ 1]^in[94];//2 inputs
        syndrom[ 3] = in[ 1]^in[95];//2 inputs
        syndrom[ 4] = in[ 2]^in[92];//2 inputs
        syndrom[ 5] = in[ 2]^in[93];//2 inputs
        syndrom[ 6] = in[ 3]^in[92];//2 inputs
        syndrom[ 7] = in[ 3]^in[93];//2 inputs
        syndrom[ 8] = in[ 4]^in[90];//2 inputs
        syndrom[ 9] = in[ 4]^in[91];//2 inputs
        syndrom[10] = in[ 5]^in[90];//2 inputs
        syndrom[11] = in[ 5]^in[91];//2 inputs
        syndrom[12] = in[ 6]^in[88];//2 inputs
        syndrom[13] = in[ 6]^in[89];//2 inputs
        syndrom[14] = in[ 7]^in[88];//2 inputs
        syndrom[15] = in[ 7]^in[89];//2 inputs
        syndrom[16] = in[ 8]^in[86];//2 inputs
        syndrom[17] = in[ 8]^in[87];//2 inputs
        syndrom[18] = in[ 9]^in[86];//2 inputs
        syndrom[19] = in[ 9]^in[87];//2 inputs
        syndrom[20] = in[10]^in[84];//2 inputs
        syndrom[21] = in[10]^in[85];//2 inputs
        syndrom[22] = in[11]^in[84];//2 inputs
        syndrom[23] = in[11]^in[85];//2 inputs
        syndrom[24] = in[12]^in[82];//2 inputs
        syndrom[25] = in[12]^in[83];//2 inputs
        syndrom[26] = in[13]^in[82];//2 inputs
        syndrom[27] = in[13]^in[83];//2 inputs
        syndrom[28] = in[14]^in[80];//2 inputs
        syndrom[29] = in[14]^in[81];//2 inputs
        syndrom[30] = in[15]^in[80];//2 inputs
        syndrom[31] = in[15]^in[81];//2 inputs
        syndrom[32] = in[16]^in[78];//2 inputs
        syndrom[33] = in[16]^in[79];//2 inputs
        syndrom[34] = in[17]^in[78];//2 inputs
        syndrom[35] = in[17]^in[79];//2 inputs
        syndrom[36] = in[18]^in[76];//2 inputs
        syndrom[37] = in[18]^in[77];//2 inputs
        syndrom[38] = in[19]^in[76];//2 inputs
        syndrom[39] = in[19]^in[77];//2 inputs
        syndrom[40] = in[20]^in[74];//2 inputs
        syndrom[41] = in[20]^in[75];//2 inputs
        syndrom[42] = in[21]^in[74];//2 inputs
        syndrom[43] = in[21]^in[75];//2 inputs
        syndrom[44] = in[22]^in[72];//2 inputs
        syndrom[45] = in[22]^in[73];//2 inputs
        syndrom[46] = in[23]^in[72];//2 inputs
        syndrom[47] = in[23]^in[73];//2 inputs
        syndrom[48] = in[24]^in[70];//2 inputs
        syndrom[49] = in[24]^in[71];//2 inputs
        syndrom[50] = in[25]^in[70];//2 inputs
        syndrom[51] = in[25]^in[71];//2 inputs
        syndrom[52] = in[26]^in[68];//2 inputs
        syndrom[53] = in[26]^in[69];//2 inputs
        syndrom[54] = in[27]^in[68];//2 inputs
        syndrom[55] = in[27]^in[69];//2 inputs
        syndrom[56] = in[28]^in[66];//2 inputs
        syndrom[57] = in[28]^in[67];//2 inputs
        syndrom[58] = in[29]^in[66];//2 inputs
        syndrom[59] = in[29]^in[67];//2 inputs
        syndrom[60] = in[30]^in[64];//2 inputs
        syndrom[61] = in[30]^in[65];//2 inputs
        syndrom[62] = in[31]^in[64];//2 inputs
        syndrom[63] = in[31]^in[65];//2 inputs
        syndrom[64] = in[32]^in[62];//2 inputs
        syndrom[65] = in[32]^in[63];//2 inputs
        syndrom[66] = in[33]^in[62];//2 inputs
        syndrom[67] = in[33]^in[63];//2 inputs
        syndrom[68] = in[34]^in[60];//2 inputs
        syndrom[69] = in[34]^in[61];//2 inputs
        syndrom[70] = in[35]^in[60];//2 inputs
        syndrom[71] = in[35]^in[61];//2 inputs
        syndrom[72] = in[36]^in[58];//2 inputs
        syndrom[73] = in[36]^in[59];//2 inputs
        syndrom[74] = in[37]^in[58];//2 inputs
        syndrom[75] = in[37]^in[59];//2 inputs
        syndrom[76] = in[38]^in[56];//2 inputs
        syndrom[77] = in[38]^in[57];//2 inputs
        syndrom[78] = in[39]^in[56];//2 inputs
        syndrom[79] = in[39]^in[57];//2 inputs
        syndrom[80] = in[40]^in[54];//2 inputs
        syndrom[81] = in[40]^in[55];//2 inputs
        syndrom[82] = in[41]^in[54];//2 inputs
        syndrom[83] = in[41]^in[55];//2 inputs
        syndrom[84] = in[42]^in[52];//2 inputs
        syndrom[85] = in[42]^in[53];//2 inputs
        syndrom[86] = in[43]^in[52];//2 inputs
        syndrom[87] = in[43]^in[53];//2 inputs
        syndrom[88] = in[44]^in[50];//2 inputs
        syndrom[89] = in[44]^in[51];//2 inputs
        syndrom[90] = in[45]^in[50];//2 inputs
        syndrom[91] = in[45]^in[51];//2 inputs
        syndrom[92] = in[46]^in[48];//2 inputs
        syndrom[93] = in[46]^in[49];//2 inputs
        syndrom[94] = in[47]^in[48];//2 inputs
        syndrom[95] = in[47]^in[49];//2 inputs
        hamming_code_192_96_f = syndrom;
    end
endfunction
wire [96-1:0] stored_data_edc = hamming_code_192_96_f(i_stored_data);
wire [96-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_96_min_delay (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [96-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [96-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_192_96_f
//Compute 96 bits Error Detection Code from a 96 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 48 49 50)
//  input bit 17 used  3 times (syndrom bits 51 52 53)
//  input bit 18 used  3 times (syndrom bits 54 55 56)
//  input bit 19 used  3 times (syndrom bits 57 58 59)
//  input bit 20 used  3 times (syndrom bits 60 61 62)
//  input bit 21 used  3 times (syndrom bits 63 64 65)
//  input bit 22 used  3 times (syndrom bits 66 67 68)
//  input bit 23 used  3 times (syndrom bits 69 70 71)
//  input bit 24 used  3 times (syndrom bits 72 73 74)
//  input bit 25 used  3 times (syndrom bits 75 76 77)
//  input bit 26 used  3 times (syndrom bits 78 79 80)
//  input bit 27 used  3 times (syndrom bits 81 82 83)
//  input bit 28 used  3 times (syndrom bits 84 85 86)
//  input bit 29 used  3 times (syndrom bits 87 88 89)
//  input bit 30 used  3 times (syndrom bits 90 91 92)
//  input bit 31 used  3 times (syndrom bits 93 94 95)
//  input bit 32 used  3 times (syndrom bits 90 93 94)
//  input bit 33 used  3 times (syndrom bits 91 92 95)
//  input bit 34 used  3 times (syndrom bits 84 87 88)
//  input bit 35 used  3 times (syndrom bits 85 86 89)
//  input bit 36 used  3 times (syndrom bits 78 81 82)
//  input bit 37 used  3 times (syndrom bits 79 80 83)
//  input bit 38 used  3 times (syndrom bits 72 75 76)
//  input bit 39 used  3 times (syndrom bits 73 74 77)
//  input bit 40 used  3 times (syndrom bits 66 69 70)
//  input bit 41 used  3 times (syndrom bits 67 68 71)
//  input bit 42 used  3 times (syndrom bits 60 63 64)
//  input bit 43 used  3 times (syndrom bits 61 62 65)
//  input bit 44 used  3 times (syndrom bits 54 57 58)
//  input bit 45 used  3 times (syndrom bits 55 56 59)
//  input bit 46 used  3 times (syndrom bits 48 51 52)
//  input bit 47 used  3 times (syndrom bits 49 50 53)
//  input bit 48 used  3 times (syndrom bits 42 45 46)
//  input bit 49 used  3 times (syndrom bits 43 44 47)
//  input bit 50 used  3 times (syndrom bits 36 39 40)
//  input bit 51 used  3 times (syndrom bits 37 38 41)
//  input bit 52 used  3 times (syndrom bits 30 33 34)
//  input bit 53 used  3 times (syndrom bits 31 32 35)
//  input bit 54 used  3 times (syndrom bits 24 27 28)
//  input bit 55 used  3 times (syndrom bits 25 26 29)
//  input bit 56 used  3 times (syndrom bits 18 21 22)
//  input bit 57 used  3 times (syndrom bits 19 20 23)
//  input bit 58 used  3 times (syndrom bits 12 15 16)
//  input bit 59 used  3 times (syndrom bits 13 14 17)
//  input bit 60 used  3 times (syndrom bits 6 9 10)
//  input bit 61 used  3 times (syndrom bits 7 8 11)
//  input bit 62 used  3 times (syndrom bits 0 3 4)
//  input bit 63 used  3 times (syndrom bits 1 2 5)
//  input bit 64 used  3 times (syndrom bits 1 3 5)
//  input bit 65 used  3 times (syndrom bits 0 2 4)
//  input bit 66 used  3 times (syndrom bits 7 9 11)
//  input bit 67 used  3 times (syndrom bits 6 8 10)
//  input bit 68 used  3 times (syndrom bits 13 15 17)
//  input bit 69 used  3 times (syndrom bits 12 14 16)
//  input bit 70 used  3 times (syndrom bits 19 21 23)
//  input bit 71 used  3 times (syndrom bits 18 20 22)
//  input bit 72 used  3 times (syndrom bits 25 27 29)
//  input bit 73 used  3 times (syndrom bits 24 26 28)
//  input bit 74 used  3 times (syndrom bits 31 33 35)
//  input bit 75 used  3 times (syndrom bits 30 32 34)
//  input bit 76 used  3 times (syndrom bits 37 39 41)
//  input bit 77 used  3 times (syndrom bits 36 38 40)
//  input bit 78 used  3 times (syndrom bits 43 45 47)
//  input bit 79 used  3 times (syndrom bits 42 44 46)
//  input bit 80 used  3 times (syndrom bits 49 51 53)
//  input bit 81 used  3 times (syndrom bits 48 50 52)
//  input bit 82 used  3 times (syndrom bits 55 57 59)
//  input bit 83 used  3 times (syndrom bits 54 56 58)
//  input bit 84 used  3 times (syndrom bits 61 63 65)
//  input bit 85 used  3 times (syndrom bits 60 62 64)
//  input bit 86 used  3 times (syndrom bits 67 69 71)
//  input bit 87 used  3 times (syndrom bits 66 68 70)
//  input bit 88 used  3 times (syndrom bits 73 75 77)
//  input bit 89 used  3 times (syndrom bits 72 74 76)
//  input bit 90 used  3 times (syndrom bits 79 81 83)
//  input bit 91 used  3 times (syndrom bits 78 80 82)
//  input bit 92 used  3 times (syndrom bits 85 87 89)
//  input bit 93 used  3 times (syndrom bits 84 86 88)
//  input bit 94 used  3 times (syndrom bits 91 93 95)
//  input bit 95 used  3 times (syndrom bits 90 92 94)
function [96-1:0] extended_hamming_code_192_96_f;
    input [96-1:0] in;
    reg [96-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[62]^in[65];//3 inputs
        syndrom[ 1] = in[ 0]^in[63]^in[64];//3 inputs
        syndrom[ 2] = in[ 0]^in[63]^in[65];//3 inputs
        syndrom[ 3] = in[ 1]^in[62]^in[64];//3 inputs
        syndrom[ 4] = in[ 1]^in[62]^in[65];//3 inputs
        syndrom[ 5] = in[ 1]^in[63]^in[64];//3 inputs
        syndrom[ 6] = in[ 2]^in[60]^in[67];//3 inputs
        syndrom[ 7] = in[ 2]^in[61]^in[66];//3 inputs
        syndrom[ 8] = in[ 2]^in[61]^in[67];//3 inputs
        syndrom[ 9] = in[ 3]^in[60]^in[66];//3 inputs
        syndrom[10] = in[ 3]^in[60]^in[67];//3 inputs
        syndrom[11] = in[ 3]^in[61]^in[66];//3 inputs
        syndrom[12] = in[ 4]^in[58]^in[69];//3 inputs
        syndrom[13] = in[ 4]^in[59]^in[68];//3 inputs
        syndrom[14] = in[ 4]^in[59]^in[69];//3 inputs
        syndrom[15] = in[ 5]^in[58]^in[68];//3 inputs
        syndrom[16] = in[ 5]^in[58]^in[69];//3 inputs
        syndrom[17] = in[ 5]^in[59]^in[68];//3 inputs
        syndrom[18] = in[ 6]^in[56]^in[71];//3 inputs
        syndrom[19] = in[ 6]^in[57]^in[70];//3 inputs
        syndrom[20] = in[ 6]^in[57]^in[71];//3 inputs
        syndrom[21] = in[ 7]^in[56]^in[70];//3 inputs
        syndrom[22] = in[ 7]^in[56]^in[71];//3 inputs
        syndrom[23] = in[ 7]^in[57]^in[70];//3 inputs
        syndrom[24] = in[ 8]^in[54]^in[73];//3 inputs
        syndrom[25] = in[ 8]^in[55]^in[72];//3 inputs
        syndrom[26] = in[ 8]^in[55]^in[73];//3 inputs
        syndrom[27] = in[ 9]^in[54]^in[72];//3 inputs
        syndrom[28] = in[ 9]^in[54]^in[73];//3 inputs
        syndrom[29] = in[ 9]^in[55]^in[72];//3 inputs
        syndrom[30] = in[10]^in[52]^in[75];//3 inputs
        syndrom[31] = in[10]^in[53]^in[74];//3 inputs
        syndrom[32] = in[10]^in[53]^in[75];//3 inputs
        syndrom[33] = in[11]^in[52]^in[74];//3 inputs
        syndrom[34] = in[11]^in[52]^in[75];//3 inputs
        syndrom[35] = in[11]^in[53]^in[74];//3 inputs
        syndrom[36] = in[12]^in[50]^in[77];//3 inputs
        syndrom[37] = in[12]^in[51]^in[76];//3 inputs
        syndrom[38] = in[12]^in[51]^in[77];//3 inputs
        syndrom[39] = in[13]^in[50]^in[76];//3 inputs
        syndrom[40] = in[13]^in[50]^in[77];//3 inputs
        syndrom[41] = in[13]^in[51]^in[76];//3 inputs
        syndrom[42] = in[14]^in[48]^in[79];//3 inputs
        syndrom[43] = in[14]^in[49]^in[78];//3 inputs
        syndrom[44] = in[14]^in[49]^in[79];//3 inputs
        syndrom[45] = in[15]^in[48]^in[78];//3 inputs
        syndrom[46] = in[15]^in[48]^in[79];//3 inputs
        syndrom[47] = in[15]^in[49]^in[78];//3 inputs
        syndrom[48] = in[16]^in[46]^in[81];//3 inputs
        syndrom[49] = in[16]^in[47]^in[80];//3 inputs
        syndrom[50] = in[16]^in[47]^in[81];//3 inputs
        syndrom[51] = in[17]^in[46]^in[80];//3 inputs
        syndrom[52] = in[17]^in[46]^in[81];//3 inputs
        syndrom[53] = in[17]^in[47]^in[80];//3 inputs
        syndrom[54] = in[18]^in[44]^in[83];//3 inputs
        syndrom[55] = in[18]^in[45]^in[82];//3 inputs
        syndrom[56] = in[18]^in[45]^in[83];//3 inputs
        syndrom[57] = in[19]^in[44]^in[82];//3 inputs
        syndrom[58] = in[19]^in[44]^in[83];//3 inputs
        syndrom[59] = in[19]^in[45]^in[82];//3 inputs
        syndrom[60] = in[20]^in[42]^in[85];//3 inputs
        syndrom[61] = in[20]^in[43]^in[84];//3 inputs
        syndrom[62] = in[20]^in[43]^in[85];//3 inputs
        syndrom[63] = in[21]^in[42]^in[84];//3 inputs
        syndrom[64] = in[21]^in[42]^in[85];//3 inputs
        syndrom[65] = in[21]^in[43]^in[84];//3 inputs
        syndrom[66] = in[22]^in[40]^in[87];//3 inputs
        syndrom[67] = in[22]^in[41]^in[86];//3 inputs
        syndrom[68] = in[22]^in[41]^in[87];//3 inputs
        syndrom[69] = in[23]^in[40]^in[86];//3 inputs
        syndrom[70] = in[23]^in[40]^in[87];//3 inputs
        syndrom[71] = in[23]^in[41]^in[86];//3 inputs
        syndrom[72] = in[24]^in[38]^in[89];//3 inputs
        syndrom[73] = in[24]^in[39]^in[88];//3 inputs
        syndrom[74] = in[24]^in[39]^in[89];//3 inputs
        syndrom[75] = in[25]^in[38]^in[88];//3 inputs
        syndrom[76] = in[25]^in[38]^in[89];//3 inputs
        syndrom[77] = in[25]^in[39]^in[88];//3 inputs
        syndrom[78] = in[26]^in[36]^in[91];//3 inputs
        syndrom[79] = in[26]^in[37]^in[90];//3 inputs
        syndrom[80] = in[26]^in[37]^in[91];//3 inputs
        syndrom[81] = in[27]^in[36]^in[90];//3 inputs
        syndrom[82] = in[27]^in[36]^in[91];//3 inputs
        syndrom[83] = in[27]^in[37]^in[90];//3 inputs
        syndrom[84] = in[28]^in[34]^in[93];//3 inputs
        syndrom[85] = in[28]^in[35]^in[92];//3 inputs
        syndrom[86] = in[28]^in[35]^in[93];//3 inputs
        syndrom[87] = in[29]^in[34]^in[92];//3 inputs
        syndrom[88] = in[29]^in[34]^in[93];//3 inputs
        syndrom[89] = in[29]^in[35]^in[92];//3 inputs
        syndrom[90] = in[30]^in[32]^in[95];//3 inputs
        syndrom[91] = in[30]^in[33]^in[94];//3 inputs
        syndrom[92] = in[30]^in[33]^in[95];//3 inputs
        syndrom[93] = in[31]^in[32]^in[94];//3 inputs
        syndrom[94] = in[31]^in[32]^in[95];//3 inputs
        syndrom[95] = in[31]^in[33]^in[94];//3 inputs
        extended_hamming_code_192_96_f = syndrom;
    end
endfunction
wire [96-1:0] stored_data_edc = extended_hamming_code_192_96_f(i_stored_data);
wire [96-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_96_min_delay (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [96-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [96-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [96-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_192_96_f
//Compute 96 bits Error Detection Code from a 96 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 48 49 50)
//  input bit 17 used  3 times (syndrom bits 51 52 53)
//  input bit 18 used  3 times (syndrom bits 54 55 56)
//  input bit 19 used  3 times (syndrom bits 57 58 59)
//  input bit 20 used  3 times (syndrom bits 60 61 62)
//  input bit 21 used  3 times (syndrom bits 63 64 65)
//  input bit 22 used  3 times (syndrom bits 66 67 68)
//  input bit 23 used  3 times (syndrom bits 69 70 71)
//  input bit 24 used  3 times (syndrom bits 72 73 74)
//  input bit 25 used  3 times (syndrom bits 75 76 77)
//  input bit 26 used  3 times (syndrom bits 78 79 80)
//  input bit 27 used  3 times (syndrom bits 81 82 83)
//  input bit 28 used  3 times (syndrom bits 84 85 86)
//  input bit 29 used  3 times (syndrom bits 87 88 89)
//  input bit 30 used  3 times (syndrom bits 90 91 92)
//  input bit 31 used  3 times (syndrom bits 93 94 95)
//  input bit 32 used  3 times (syndrom bits 90 93 94)
//  input bit 33 used  3 times (syndrom bits 91 92 95)
//  input bit 34 used  3 times (syndrom bits 84 87 88)
//  input bit 35 used  3 times (syndrom bits 85 86 89)
//  input bit 36 used  3 times (syndrom bits 78 81 82)
//  input bit 37 used  3 times (syndrom bits 79 80 83)
//  input bit 38 used  3 times (syndrom bits 72 75 76)
//  input bit 39 used  3 times (syndrom bits 73 74 77)
//  input bit 40 used  3 times (syndrom bits 66 69 70)
//  input bit 41 used  3 times (syndrom bits 67 68 71)
//  input bit 42 used  3 times (syndrom bits 60 63 64)
//  input bit 43 used  3 times (syndrom bits 61 62 65)
//  input bit 44 used  3 times (syndrom bits 54 57 58)
//  input bit 45 used  3 times (syndrom bits 55 56 59)
//  input bit 46 used  3 times (syndrom bits 48 51 52)
//  input bit 47 used  3 times (syndrom bits 49 50 53)
//  input bit 48 used  3 times (syndrom bits 42 45 46)
//  input bit 49 used  3 times (syndrom bits 43 44 47)
//  input bit 50 used  3 times (syndrom bits 36 39 40)
//  input bit 51 used  3 times (syndrom bits 37 38 41)
//  input bit 52 used  3 times (syndrom bits 30 33 34)
//  input bit 53 used  3 times (syndrom bits 31 32 35)
//  input bit 54 used  3 times (syndrom bits 24 27 28)
//  input bit 55 used  3 times (syndrom bits 25 26 29)
//  input bit 56 used  3 times (syndrom bits 18 21 22)
//  input bit 57 used  3 times (syndrom bits 19 20 23)
//  input bit 58 used  3 times (syndrom bits 12 15 16)
//  input bit 59 used  3 times (syndrom bits 13 14 17)
//  input bit 60 used  3 times (syndrom bits 6 9 10)
//  input bit 61 used  3 times (syndrom bits 7 8 11)
//  input bit 62 used  3 times (syndrom bits 0 3 4)
//  input bit 63 used  3 times (syndrom bits 1 2 5)
//  input bit 64 used  3 times (syndrom bits 1 3 5)
//  input bit 65 used  3 times (syndrom bits 0 2 4)
//  input bit 66 used  3 times (syndrom bits 7 9 11)
//  input bit 67 used  3 times (syndrom bits 6 8 10)
//  input bit 68 used  3 times (syndrom bits 13 15 17)
//  input bit 69 used  3 times (syndrom bits 12 14 16)
//  input bit 70 used  3 times (syndrom bits 19 21 23)
//  input bit 71 used  3 times (syndrom bits 18 20 22)
//  input bit 72 used  3 times (syndrom bits 25 27 29)
//  input bit 73 used  3 times (syndrom bits 24 26 28)
//  input bit 74 used  3 times (syndrom bits 31 33 35)
//  input bit 75 used  3 times (syndrom bits 30 32 34)
//  input bit 76 used  3 times (syndrom bits 37 39 41)
//  input bit 77 used  3 times (syndrom bits 36 38 40)
//  input bit 78 used  3 times (syndrom bits 43 45 47)
//  input bit 79 used  3 times (syndrom bits 42 44 46)
//  input bit 80 used  3 times (syndrom bits 49 51 53)
//  input bit 81 used  3 times (syndrom bits 48 50 52)
//  input bit 82 used  3 times (syndrom bits 55 57 59)
//  input bit 83 used  3 times (syndrom bits 54 56 58)
//  input bit 84 used  3 times (syndrom bits 61 63 65)
//  input bit 85 used  3 times (syndrom bits 60 62 64)
//  input bit 86 used  3 times (syndrom bits 67 69 71)
//  input bit 87 used  3 times (syndrom bits 66 68 70)
//  input bit 88 used  3 times (syndrom bits 73 75 77)
//  input bit 89 used  3 times (syndrom bits 72 74 76)
//  input bit 90 used  3 times (syndrom bits 79 81 83)
//  input bit 91 used  3 times (syndrom bits 78 80 82)
//  input bit 92 used  3 times (syndrom bits 85 87 89)
//  input bit 93 used  3 times (syndrom bits 84 86 88)
//  input bit 94 used  3 times (syndrom bits 91 93 95)
//  input bit 95 used  3 times (syndrom bits 90 92 94)
function [96-1:0] extended_hamming_code_192_96_f;
    input [96-1:0] in;
    reg [96-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[62]^in[65];//3 inputs
        syndrom[ 1] = in[ 0]^in[63]^in[64];//3 inputs
        syndrom[ 2] = in[ 0]^in[63]^in[65];//3 inputs
        syndrom[ 3] = in[ 1]^in[62]^in[64];//3 inputs
        syndrom[ 4] = in[ 1]^in[62]^in[65];//3 inputs
        syndrom[ 5] = in[ 1]^in[63]^in[64];//3 inputs
        syndrom[ 6] = in[ 2]^in[60]^in[67];//3 inputs
        syndrom[ 7] = in[ 2]^in[61]^in[66];//3 inputs
        syndrom[ 8] = in[ 2]^in[61]^in[67];//3 inputs
        syndrom[ 9] = in[ 3]^in[60]^in[66];//3 inputs
        syndrom[10] = in[ 3]^in[60]^in[67];//3 inputs
        syndrom[11] = in[ 3]^in[61]^in[66];//3 inputs
        syndrom[12] = in[ 4]^in[58]^in[69];//3 inputs
        syndrom[13] = in[ 4]^in[59]^in[68];//3 inputs
        syndrom[14] = in[ 4]^in[59]^in[69];//3 inputs
        syndrom[15] = in[ 5]^in[58]^in[68];//3 inputs
        syndrom[16] = in[ 5]^in[58]^in[69];//3 inputs
        syndrom[17] = in[ 5]^in[59]^in[68];//3 inputs
        syndrom[18] = in[ 6]^in[56]^in[71];//3 inputs
        syndrom[19] = in[ 6]^in[57]^in[70];//3 inputs
        syndrom[20] = in[ 6]^in[57]^in[71];//3 inputs
        syndrom[21] = in[ 7]^in[56]^in[70];//3 inputs
        syndrom[22] = in[ 7]^in[56]^in[71];//3 inputs
        syndrom[23] = in[ 7]^in[57]^in[70];//3 inputs
        syndrom[24] = in[ 8]^in[54]^in[73];//3 inputs
        syndrom[25] = in[ 8]^in[55]^in[72];//3 inputs
        syndrom[26] = in[ 8]^in[55]^in[73];//3 inputs
        syndrom[27] = in[ 9]^in[54]^in[72];//3 inputs
        syndrom[28] = in[ 9]^in[54]^in[73];//3 inputs
        syndrom[29] = in[ 9]^in[55]^in[72];//3 inputs
        syndrom[30] = in[10]^in[52]^in[75];//3 inputs
        syndrom[31] = in[10]^in[53]^in[74];//3 inputs
        syndrom[32] = in[10]^in[53]^in[75];//3 inputs
        syndrom[33] = in[11]^in[52]^in[74];//3 inputs
        syndrom[34] = in[11]^in[52]^in[75];//3 inputs
        syndrom[35] = in[11]^in[53]^in[74];//3 inputs
        syndrom[36] = in[12]^in[50]^in[77];//3 inputs
        syndrom[37] = in[12]^in[51]^in[76];//3 inputs
        syndrom[38] = in[12]^in[51]^in[77];//3 inputs
        syndrom[39] = in[13]^in[50]^in[76];//3 inputs
        syndrom[40] = in[13]^in[50]^in[77];//3 inputs
        syndrom[41] = in[13]^in[51]^in[76];//3 inputs
        syndrom[42] = in[14]^in[48]^in[79];//3 inputs
        syndrom[43] = in[14]^in[49]^in[78];//3 inputs
        syndrom[44] = in[14]^in[49]^in[79];//3 inputs
        syndrom[45] = in[15]^in[48]^in[78];//3 inputs
        syndrom[46] = in[15]^in[48]^in[79];//3 inputs
        syndrom[47] = in[15]^in[49]^in[78];//3 inputs
        syndrom[48] = in[16]^in[46]^in[81];//3 inputs
        syndrom[49] = in[16]^in[47]^in[80];//3 inputs
        syndrom[50] = in[16]^in[47]^in[81];//3 inputs
        syndrom[51] = in[17]^in[46]^in[80];//3 inputs
        syndrom[52] = in[17]^in[46]^in[81];//3 inputs
        syndrom[53] = in[17]^in[47]^in[80];//3 inputs
        syndrom[54] = in[18]^in[44]^in[83];//3 inputs
        syndrom[55] = in[18]^in[45]^in[82];//3 inputs
        syndrom[56] = in[18]^in[45]^in[83];//3 inputs
        syndrom[57] = in[19]^in[44]^in[82];//3 inputs
        syndrom[58] = in[19]^in[44]^in[83];//3 inputs
        syndrom[59] = in[19]^in[45]^in[82];//3 inputs
        syndrom[60] = in[20]^in[42]^in[85];//3 inputs
        syndrom[61] = in[20]^in[43]^in[84];//3 inputs
        syndrom[62] = in[20]^in[43]^in[85];//3 inputs
        syndrom[63] = in[21]^in[42]^in[84];//3 inputs
        syndrom[64] = in[21]^in[42]^in[85];//3 inputs
        syndrom[65] = in[21]^in[43]^in[84];//3 inputs
        syndrom[66] = in[22]^in[40]^in[87];//3 inputs
        syndrom[67] = in[22]^in[41]^in[86];//3 inputs
        syndrom[68] = in[22]^in[41]^in[87];//3 inputs
        syndrom[69] = in[23]^in[40]^in[86];//3 inputs
        syndrom[70] = in[23]^in[40]^in[87];//3 inputs
        syndrom[71] = in[23]^in[41]^in[86];//3 inputs
        syndrom[72] = in[24]^in[38]^in[89];//3 inputs
        syndrom[73] = in[24]^in[39]^in[88];//3 inputs
        syndrom[74] = in[24]^in[39]^in[89];//3 inputs
        syndrom[75] = in[25]^in[38]^in[88];//3 inputs
        syndrom[76] = in[25]^in[38]^in[89];//3 inputs
        syndrom[77] = in[25]^in[39]^in[88];//3 inputs
        syndrom[78] = in[26]^in[36]^in[91];//3 inputs
        syndrom[79] = in[26]^in[37]^in[90];//3 inputs
        syndrom[80] = in[26]^in[37]^in[91];//3 inputs
        syndrom[81] = in[27]^in[36]^in[90];//3 inputs
        syndrom[82] = in[27]^in[36]^in[91];//3 inputs
        syndrom[83] = in[27]^in[37]^in[90];//3 inputs
        syndrom[84] = in[28]^in[34]^in[93];//3 inputs
        syndrom[85] = in[28]^in[35]^in[92];//3 inputs
        syndrom[86] = in[28]^in[35]^in[93];//3 inputs
        syndrom[87] = in[29]^in[34]^in[92];//3 inputs
        syndrom[88] = in[29]^in[34]^in[93];//3 inputs
        syndrom[89] = in[29]^in[35]^in[92];//3 inputs
        syndrom[90] = in[30]^in[32]^in[95];//3 inputs
        syndrom[91] = in[30]^in[33]^in[94];//3 inputs
        syndrom[92] = in[30]^in[33]^in[95];//3 inputs
        syndrom[93] = in[31]^in[32]^in[94];//3 inputs
        syndrom[94] = in[31]^in[32]^in[95];//3 inputs
        syndrom[95] = in[31]^in[33]^in[94];//3 inputs
        extended_hamming_code_192_96_f = syndrom;
    end
endfunction
function [2+96-1:0] extended_hamming_code_192_96_f_correction_pattern_f;
    input [96-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [96-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {96{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {96{1'b0}};
			end	
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 0]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 1]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 2]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 3]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 4]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 5]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 6]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 7]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 8]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 9]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[10]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[11]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[12]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[13]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[14]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[15]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[16]=1'b1;
			end
			96'b000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[17]=1'b1;
			end
			96'b000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[18]=1'b1;
			end
			96'b000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[19]=1'b1;
			end
			96'b000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[20]=1'b1;
			end
			96'b000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[21]=1'b1;
			end
			96'b000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[22]=1'b1;
			end
			96'b000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[23]=1'b1;
			end
			96'b000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[24]=1'b1;
			end
			96'b000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[25]=1'b1;
			end
			96'b000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[26]=1'b1;
			end
			96'b000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[27]=1'b1;
			end
			96'b000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[28]=1'b1;
			end
			96'b000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[29]=1'b1;
			end
			96'b000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[30]=1'b1;
			end
			96'b111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[31]=1'b1;
			end
			96'b011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[32]=1'b1;
			end
			96'b100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[33]=1'b1;
			end
			96'b000000011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[34]=1'b1;
			end
			96'b000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[35]=1'b1;
			end
			96'b000000000000011001000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[36]=1'b1;
			end
			96'b000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[37]=1'b1;
			end
			96'b000000000000000000011001000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[38]=1'b1;
			end
			96'b000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[39]=1'b1;
			end
			96'b000000000000000000000000011001000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[40]=1'b1;
			end
			96'b000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[41]=1'b1;
			end
			96'b000000000000000000000000000000011001000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[42]=1'b1;
			end
			96'b000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[43]=1'b1;
			end
			96'b000000000000000000000000000000000000011001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[44]=1'b1;
			end
			96'b000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[45]=1'b1;
			end
			96'b000000000000000000000000000000000000000000011001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[46]=1'b1;
			end
			96'b000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[47]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000011001000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[48]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[49]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000011001000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[50]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[51]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000011001000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[52]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[53]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000011001000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[54]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000100110000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[55]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000011001000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[56]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000100110000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[57]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[58]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[59]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[60]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[61]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001: begin
				correction_pattern = {96{1'b0}};correction_pattern[62]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110: begin
				correction_pattern = {96{1'b0}};correction_pattern[63]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010: begin
				correction_pattern = {96{1'b0}};correction_pattern[64]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101: begin
				correction_pattern = {96{1'b0}};correction_pattern[65]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[66]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[67]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[68]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[69]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[70]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000010101000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[71]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[72]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000010101000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[73]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[74]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000010101000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[75]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[76]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000010101000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[77]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[78]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000010101000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[79]=1'b1;
			end
			96'b000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[80]=1'b1;
			end
			96'b000000000000000000000000000000000000000000010101000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[81]=1'b1;
			end
			96'b000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[82]=1'b1;
			end
			96'b000000000000000000000000000000000000010101000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[83]=1'b1;
			end
			96'b000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[84]=1'b1;
			end
			96'b000000000000000000000000000000010101000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[85]=1'b1;
			end
			96'b000000000000000000000000101010000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[86]=1'b1;
			end
			96'b000000000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[87]=1'b1;
			end
			96'b000000000000000000101010000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[88]=1'b1;
			end
			96'b000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[89]=1'b1;
			end
			96'b000000000000101010000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[90]=1'b1;
			end
			96'b000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[91]=1'b1;
			end
			96'b000000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[92]=1'b1;
			end
			96'b000000010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[93]=1'b1;
			end
			96'b101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[94]=1'b1;
			end
			96'b010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[95]=1'b1;
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			96'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_192_96_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [96-1:0] stored_data_edc = extended_hamming_code_192_96_f(i_stored_data);
wire [96-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [96-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_192_96_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_128_min_delay (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [128-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [128-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_256_128_f
//Compute 128 bits Error Detection Code from a 128 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used   2 times (syndrom bits 0 1)
//  input bit   1 used   2 times (syndrom bits 2 3)
//  input bit   2 used   2 times (syndrom bits 4 5)
//  input bit   3 used   2 times (syndrom bits 6 7)
//  input bit   4 used   2 times (syndrom bits 8 9)
//  input bit   5 used   2 times (syndrom bits 10 11)
//  input bit   6 used   2 times (syndrom bits 12 13)
//  input bit   7 used   2 times (syndrom bits 14 15)
//  input bit   8 used   2 times (syndrom bits 16 17)
//  input bit   9 used   2 times (syndrom bits 18 19)
//  input bit  10 used   2 times (syndrom bits 20 21)
//  input bit  11 used   2 times (syndrom bits 22 23)
//  input bit  12 used   2 times (syndrom bits 24 25)
//  input bit  13 used   2 times (syndrom bits 26 27)
//  input bit  14 used   2 times (syndrom bits 28 29)
//  input bit  15 used   2 times (syndrom bits 30 31)
//  input bit  16 used   2 times (syndrom bits 32 33)
//  input bit  17 used   2 times (syndrom bits 34 35)
//  input bit  18 used   2 times (syndrom bits 36 37)
//  input bit  19 used   2 times (syndrom bits 38 39)
//  input bit  20 used   2 times (syndrom bits 40 41)
//  input bit  21 used   2 times (syndrom bits 42 43)
//  input bit  22 used   2 times (syndrom bits 44 45)
//  input bit  23 used   2 times (syndrom bits 46 47)
//  input bit  24 used   2 times (syndrom bits 48 49)
//  input bit  25 used   2 times (syndrom bits 50 51)
//  input bit  26 used   2 times (syndrom bits 52 53)
//  input bit  27 used   2 times (syndrom bits 54 55)
//  input bit  28 used   2 times (syndrom bits 56 57)
//  input bit  29 used   2 times (syndrom bits 58 59)
//  input bit  30 used   2 times (syndrom bits 60 61)
//  input bit  31 used   2 times (syndrom bits 62 63)
//  input bit  32 used   2 times (syndrom bits 64 65)
//  input bit  33 used   2 times (syndrom bits 66 67)
//  input bit  34 used   2 times (syndrom bits 68 69)
//  input bit  35 used   2 times (syndrom bits 70 71)
//  input bit  36 used   2 times (syndrom bits 72 73)
//  input bit  37 used   2 times (syndrom bits 74 75)
//  input bit  38 used   2 times (syndrom bits 76 77)
//  input bit  39 used   2 times (syndrom bits 78 79)
//  input bit  40 used   2 times (syndrom bits 80 81)
//  input bit  41 used   2 times (syndrom bits 82 83)
//  input bit  42 used   2 times (syndrom bits 84 85)
//  input bit  43 used   2 times (syndrom bits 86 87)
//  input bit  44 used   2 times (syndrom bits 88 89)
//  input bit  45 used   2 times (syndrom bits 90 91)
//  input bit  46 used   2 times (syndrom bits 92 93)
//  input bit  47 used   2 times (syndrom bits 94 95)
//  input bit  48 used   2 times (syndrom bits 96 97)
//  input bit  49 used   2 times (syndrom bits 98 99)
//  input bit  50 used   2 times (syndrom bits 100 101)
//  input bit  51 used   2 times (syndrom bits 102 103)
//  input bit  52 used   2 times (syndrom bits 104 105)
//  input bit  53 used   2 times (syndrom bits 106 107)
//  input bit  54 used   2 times (syndrom bits 108 109)
//  input bit  55 used   2 times (syndrom bits 110 111)
//  input bit  56 used   2 times (syndrom bits 112 113)
//  input bit  57 used   2 times (syndrom bits 114 115)
//  input bit  58 used   2 times (syndrom bits 116 117)
//  input bit  59 used   2 times (syndrom bits 118 119)
//  input bit  60 used   2 times (syndrom bits 120 121)
//  input bit  61 used   2 times (syndrom bits 122 123)
//  input bit  62 used   2 times (syndrom bits 124 125)
//  input bit  63 used   2 times (syndrom bits 126 127)
//  input bit  64 used   2 times (syndrom bits 124 126)
//  input bit  65 used   2 times (syndrom bits 125 127)
//  input bit  66 used   2 times (syndrom bits 120 122)
//  input bit  67 used   2 times (syndrom bits 121 123)
//  input bit  68 used   2 times (syndrom bits 116 118)
//  input bit  69 used   2 times (syndrom bits 117 119)
//  input bit  70 used   2 times (syndrom bits 112 114)
//  input bit  71 used   2 times (syndrom bits 113 115)
//  input bit  72 used   2 times (syndrom bits 108 110)
//  input bit  73 used   2 times (syndrom bits 109 111)
//  input bit  74 used   2 times (syndrom bits 104 106)
//  input bit  75 used   2 times (syndrom bits 105 107)
//  input bit  76 used   2 times (syndrom bits 100 102)
//  input bit  77 used   2 times (syndrom bits 101 103)
//  input bit  78 used   2 times (syndrom bits 96 98)
//  input bit  79 used   2 times (syndrom bits 97 99)
//  input bit  80 used   2 times (syndrom bits 92 94)
//  input bit  81 used   2 times (syndrom bits 93 95)
//  input bit  82 used   2 times (syndrom bits 88 90)
//  input bit  83 used   2 times (syndrom bits 89 91)
//  input bit  84 used   2 times (syndrom bits 84 86)
//  input bit  85 used   2 times (syndrom bits 85 87)
//  input bit  86 used   2 times (syndrom bits 80 82)
//  input bit  87 used   2 times (syndrom bits 81 83)
//  input bit  88 used   2 times (syndrom bits 76 78)
//  input bit  89 used   2 times (syndrom bits 77 79)
//  input bit  90 used   2 times (syndrom bits 72 74)
//  input bit  91 used   2 times (syndrom bits 73 75)
//  input bit  92 used   2 times (syndrom bits 68 70)
//  input bit  93 used   2 times (syndrom bits 69 71)
//  input bit  94 used   2 times (syndrom bits 64 66)
//  input bit  95 used   2 times (syndrom bits 65 67)
//  input bit  96 used   2 times (syndrom bits 60 62)
//  input bit  97 used   2 times (syndrom bits 61 63)
//  input bit  98 used   2 times (syndrom bits 56 58)
//  input bit  99 used   2 times (syndrom bits 57 59)
//  input bit 100 used   2 times (syndrom bits 52 54)
//  input bit 101 used   2 times (syndrom bits 53 55)
//  input bit 102 used   2 times (syndrom bits 48 50)
//  input bit 103 used   2 times (syndrom bits 49 51)
//  input bit 104 used   2 times (syndrom bits 44 46)
//  input bit 105 used   2 times (syndrom bits 45 47)
//  input bit 106 used   2 times (syndrom bits 40 42)
//  input bit 107 used   2 times (syndrom bits 41 43)
//  input bit 108 used   2 times (syndrom bits 36 38)
//  input bit 109 used   2 times (syndrom bits 37 39)
//  input bit 110 used   2 times (syndrom bits 32 34)
//  input bit 111 used   2 times (syndrom bits 33 35)
//  input bit 112 used   2 times (syndrom bits 28 30)
//  input bit 113 used   2 times (syndrom bits 29 31)
//  input bit 114 used   2 times (syndrom bits 24 26)
//  input bit 115 used   2 times (syndrom bits 25 27)
//  input bit 116 used   2 times (syndrom bits 20 22)
//  input bit 117 used   2 times (syndrom bits 21 23)
//  input bit 118 used   2 times (syndrom bits 16 18)
//  input bit 119 used   2 times (syndrom bits 17 19)
//  input bit 120 used   2 times (syndrom bits 12 14)
//  input bit 121 used   2 times (syndrom bits 13 15)
//  input bit 122 used   2 times (syndrom bits 8 10)
//  input bit 123 used   2 times (syndrom bits 9 11)
//  input bit 124 used   2 times (syndrom bits 4 6)
//  input bit 125 used   2 times (syndrom bits 5 7)
//  input bit 126 used   2 times (syndrom bits 0 2)
//  input bit 127 used   2 times (syndrom bits 1 3)
function [128-1:0] hamming_code_256_128_f;
    input [128-1:0] in;
    reg [128-1:0] syndrom;
    begin
        syndrom[  0] = in[  0]^in[126];//2 inputs
        syndrom[  1] = in[  0]^in[127];//2 inputs
        syndrom[  2] = in[  1]^in[126];//2 inputs
        syndrom[  3] = in[  1]^in[127];//2 inputs
        syndrom[  4] = in[  2]^in[124];//2 inputs
        syndrom[  5] = in[  2]^in[125];//2 inputs
        syndrom[  6] = in[  3]^in[124];//2 inputs
        syndrom[  7] = in[  3]^in[125];//2 inputs
        syndrom[  8] = in[  4]^in[122];//2 inputs
        syndrom[  9] = in[  4]^in[123];//2 inputs
        syndrom[ 10] = in[  5]^in[122];//2 inputs
        syndrom[ 11] = in[  5]^in[123];//2 inputs
        syndrom[ 12] = in[  6]^in[120];//2 inputs
        syndrom[ 13] = in[  6]^in[121];//2 inputs
        syndrom[ 14] = in[  7]^in[120];//2 inputs
        syndrom[ 15] = in[  7]^in[121];//2 inputs
        syndrom[ 16] = in[  8]^in[118];//2 inputs
        syndrom[ 17] = in[  8]^in[119];//2 inputs
        syndrom[ 18] = in[  9]^in[118];//2 inputs
        syndrom[ 19] = in[  9]^in[119];//2 inputs
        syndrom[ 20] = in[ 10]^in[116];//2 inputs
        syndrom[ 21] = in[ 10]^in[117];//2 inputs
        syndrom[ 22] = in[ 11]^in[116];//2 inputs
        syndrom[ 23] = in[ 11]^in[117];//2 inputs
        syndrom[ 24] = in[ 12]^in[114];//2 inputs
        syndrom[ 25] = in[ 12]^in[115];//2 inputs
        syndrom[ 26] = in[ 13]^in[114];//2 inputs
        syndrom[ 27] = in[ 13]^in[115];//2 inputs
        syndrom[ 28] = in[ 14]^in[112];//2 inputs
        syndrom[ 29] = in[ 14]^in[113];//2 inputs
        syndrom[ 30] = in[ 15]^in[112];//2 inputs
        syndrom[ 31] = in[ 15]^in[113];//2 inputs
        syndrom[ 32] = in[ 16]^in[110];//2 inputs
        syndrom[ 33] = in[ 16]^in[111];//2 inputs
        syndrom[ 34] = in[ 17]^in[110];//2 inputs
        syndrom[ 35] = in[ 17]^in[111];//2 inputs
        syndrom[ 36] = in[ 18]^in[108];//2 inputs
        syndrom[ 37] = in[ 18]^in[109];//2 inputs
        syndrom[ 38] = in[ 19]^in[108];//2 inputs
        syndrom[ 39] = in[ 19]^in[109];//2 inputs
        syndrom[ 40] = in[ 20]^in[106];//2 inputs
        syndrom[ 41] = in[ 20]^in[107];//2 inputs
        syndrom[ 42] = in[ 21]^in[106];//2 inputs
        syndrom[ 43] = in[ 21]^in[107];//2 inputs
        syndrom[ 44] = in[ 22]^in[104];//2 inputs
        syndrom[ 45] = in[ 22]^in[105];//2 inputs
        syndrom[ 46] = in[ 23]^in[104];//2 inputs
        syndrom[ 47] = in[ 23]^in[105];//2 inputs
        syndrom[ 48] = in[ 24]^in[102];//2 inputs
        syndrom[ 49] = in[ 24]^in[103];//2 inputs
        syndrom[ 50] = in[ 25]^in[102];//2 inputs
        syndrom[ 51] = in[ 25]^in[103];//2 inputs
        syndrom[ 52] = in[ 26]^in[100];//2 inputs
        syndrom[ 53] = in[ 26]^in[101];//2 inputs
        syndrom[ 54] = in[ 27]^in[100];//2 inputs
        syndrom[ 55] = in[ 27]^in[101];//2 inputs
        syndrom[ 56] = in[ 28]^in[ 98];//2 inputs
        syndrom[ 57] = in[ 28]^in[ 99];//2 inputs
        syndrom[ 58] = in[ 29]^in[ 98];//2 inputs
        syndrom[ 59] = in[ 29]^in[ 99];//2 inputs
        syndrom[ 60] = in[ 30]^in[ 96];//2 inputs
        syndrom[ 61] = in[ 30]^in[ 97];//2 inputs
        syndrom[ 62] = in[ 31]^in[ 96];//2 inputs
        syndrom[ 63] = in[ 31]^in[ 97];//2 inputs
        syndrom[ 64] = in[ 32]^in[ 94];//2 inputs
        syndrom[ 65] = in[ 32]^in[ 95];//2 inputs
        syndrom[ 66] = in[ 33]^in[ 94];//2 inputs
        syndrom[ 67] = in[ 33]^in[ 95];//2 inputs
        syndrom[ 68] = in[ 34]^in[ 92];//2 inputs
        syndrom[ 69] = in[ 34]^in[ 93];//2 inputs
        syndrom[ 70] = in[ 35]^in[ 92];//2 inputs
        syndrom[ 71] = in[ 35]^in[ 93];//2 inputs
        syndrom[ 72] = in[ 36]^in[ 90];//2 inputs
        syndrom[ 73] = in[ 36]^in[ 91];//2 inputs
        syndrom[ 74] = in[ 37]^in[ 90];//2 inputs
        syndrom[ 75] = in[ 37]^in[ 91];//2 inputs
        syndrom[ 76] = in[ 38]^in[ 88];//2 inputs
        syndrom[ 77] = in[ 38]^in[ 89];//2 inputs
        syndrom[ 78] = in[ 39]^in[ 88];//2 inputs
        syndrom[ 79] = in[ 39]^in[ 89];//2 inputs
        syndrom[ 80] = in[ 40]^in[ 86];//2 inputs
        syndrom[ 81] = in[ 40]^in[ 87];//2 inputs
        syndrom[ 82] = in[ 41]^in[ 86];//2 inputs
        syndrom[ 83] = in[ 41]^in[ 87];//2 inputs
        syndrom[ 84] = in[ 42]^in[ 84];//2 inputs
        syndrom[ 85] = in[ 42]^in[ 85];//2 inputs
        syndrom[ 86] = in[ 43]^in[ 84];//2 inputs
        syndrom[ 87] = in[ 43]^in[ 85];//2 inputs
        syndrom[ 88] = in[ 44]^in[ 82];//2 inputs
        syndrom[ 89] = in[ 44]^in[ 83];//2 inputs
        syndrom[ 90] = in[ 45]^in[ 82];//2 inputs
        syndrom[ 91] = in[ 45]^in[ 83];//2 inputs
        syndrom[ 92] = in[ 46]^in[ 80];//2 inputs
        syndrom[ 93] = in[ 46]^in[ 81];//2 inputs
        syndrom[ 94] = in[ 47]^in[ 80];//2 inputs
        syndrom[ 95] = in[ 47]^in[ 81];//2 inputs
        syndrom[ 96] = in[ 48]^in[ 78];//2 inputs
        syndrom[ 97] = in[ 48]^in[ 79];//2 inputs
        syndrom[ 98] = in[ 49]^in[ 78];//2 inputs
        syndrom[ 99] = in[ 49]^in[ 79];//2 inputs
        syndrom[100] = in[ 50]^in[ 76];//2 inputs
        syndrom[101] = in[ 50]^in[ 77];//2 inputs
        syndrom[102] = in[ 51]^in[ 76];//2 inputs
        syndrom[103] = in[ 51]^in[ 77];//2 inputs
        syndrom[104] = in[ 52]^in[ 74];//2 inputs
        syndrom[105] = in[ 52]^in[ 75];//2 inputs
        syndrom[106] = in[ 53]^in[ 74];//2 inputs
        syndrom[107] = in[ 53]^in[ 75];//2 inputs
        syndrom[108] = in[ 54]^in[ 72];//2 inputs
        syndrom[109] = in[ 54]^in[ 73];//2 inputs
        syndrom[110] = in[ 55]^in[ 72];//2 inputs
        syndrom[111] = in[ 55]^in[ 73];//2 inputs
        syndrom[112] = in[ 56]^in[ 70];//2 inputs
        syndrom[113] = in[ 56]^in[ 71];//2 inputs
        syndrom[114] = in[ 57]^in[ 70];//2 inputs
        syndrom[115] = in[ 57]^in[ 71];//2 inputs
        syndrom[116] = in[ 58]^in[ 68];//2 inputs
        syndrom[117] = in[ 58]^in[ 69];//2 inputs
        syndrom[118] = in[ 59]^in[ 68];//2 inputs
        syndrom[119] = in[ 59]^in[ 69];//2 inputs
        syndrom[120] = in[ 60]^in[ 66];//2 inputs
        syndrom[121] = in[ 60]^in[ 67];//2 inputs
        syndrom[122] = in[ 61]^in[ 66];//2 inputs
        syndrom[123] = in[ 61]^in[ 67];//2 inputs
        syndrom[124] = in[ 62]^in[ 64];//2 inputs
        syndrom[125] = in[ 62]^in[ 65];//2 inputs
        syndrom[126] = in[ 63]^in[ 64];//2 inputs
        syndrom[127] = in[ 63]^in[ 65];//2 inputs
        hamming_code_256_128_f = syndrom;
    end
endfunction
wire [128-1:0] stored_data_edc = hamming_code_256_128_f(i_stored_data);
wire [128-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_128_min_delay (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [128-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [128-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_256_128_f
//Compute 128 bits Error Detection Code from a 128 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used   3 times (syndrom bits 0 1 2)
//  input bit   1 used   3 times (syndrom bits 3 4 5)
//  input bit   2 used   3 times (syndrom bits 6 7 8)
//  input bit   3 used   3 times (syndrom bits 9 10 11)
//  input bit   4 used   3 times (syndrom bits 12 13 14)
//  input bit   5 used   3 times (syndrom bits 15 16 17)
//  input bit   6 used   3 times (syndrom bits 18 19 20)
//  input bit   7 used   3 times (syndrom bits 21 22 23)
//  input bit   8 used   3 times (syndrom bits 24 25 26)
//  input bit   9 used   3 times (syndrom bits 27 28 29)
//  input bit  10 used   3 times (syndrom bits 30 31 32)
//  input bit  11 used   3 times (syndrom bits 33 34 35)
//  input bit  12 used   3 times (syndrom bits 36 37 38)
//  input bit  13 used   3 times (syndrom bits 39 40 41)
//  input bit  14 used   3 times (syndrom bits 42 43 44)
//  input bit  15 used   3 times (syndrom bits 45 46 47)
//  input bit  16 used   3 times (syndrom bits 48 49 50)
//  input bit  17 used   3 times (syndrom bits 51 52 53)
//  input bit  18 used   3 times (syndrom bits 54 55 56)
//  input bit  19 used   3 times (syndrom bits 57 58 59)
//  input bit  20 used   3 times (syndrom bits 60 61 62)
//  input bit  21 used   3 times (syndrom bits 63 64 65)
//  input bit  22 used   3 times (syndrom bits 66 67 68)
//  input bit  23 used   3 times (syndrom bits 69 70 71)
//  input bit  24 used   3 times (syndrom bits 72 73 74)
//  input bit  25 used   3 times (syndrom bits 75 76 77)
//  input bit  26 used   3 times (syndrom bits 78 79 80)
//  input bit  27 used   3 times (syndrom bits 81 82 83)
//  input bit  28 used   3 times (syndrom bits 84 85 86)
//  input bit  29 used   3 times (syndrom bits 87 88 89)
//  input bit  30 used   3 times (syndrom bits 90 91 92)
//  input bit  31 used   3 times (syndrom bits 93 94 95)
//  input bit  32 used   3 times (syndrom bits 96 97 98)
//  input bit  33 used   3 times (syndrom bits 99 100 101)
//  input bit  34 used   3 times (syndrom bits 102 103 104)
//  input bit  35 used   3 times (syndrom bits 105 106 107)
//  input bit  36 used   3 times (syndrom bits 108 109 110)
//  input bit  37 used   3 times (syndrom bits 111 112 113)
//  input bit  38 used   3 times (syndrom bits 114 115 116)
//  input bit  39 used   3 times (syndrom bits 117 118 119)
//  input bit  40 used   3 times (syndrom bits 120 121 122)
//  input bit  41 used   3 times (syndrom bits 123 124 125)
//  input bit  42 used   3 times (syndrom bits 123 126 127)
//  input bit  43 used   3 times (syndrom bits 124 126 127)
//  input bit  44 used   3 times (syndrom bits 120 121 125)
//  input bit  45 used   3 times (syndrom bits 117 118 122)
//  input bit  46 used   3 times (syndrom bits 114 115 119)
//  input bit  47 used   3 times (syndrom bits 111 112 116)
//  input bit  48 used   3 times (syndrom bits 108 109 113)
//  input bit  49 used   3 times (syndrom bits 105 106 110)
//  input bit  50 used   3 times (syndrom bits 102 103 107)
//  input bit  51 used   3 times (syndrom bits 99 100 104)
//  input bit  52 used   3 times (syndrom bits 96 97 101)
//  input bit  53 used   3 times (syndrom bits 93 94 98)
//  input bit  54 used   3 times (syndrom bits 90 91 95)
//  input bit  55 used   3 times (syndrom bits 87 88 92)
//  input bit  56 used   3 times (syndrom bits 84 85 89)
//  input bit  57 used   3 times (syndrom bits 81 82 86)
//  input bit  58 used   3 times (syndrom bits 78 79 83)
//  input bit  59 used   3 times (syndrom bits 75 76 80)
//  input bit  60 used   3 times (syndrom bits 72 73 77)
//  input bit  61 used   3 times (syndrom bits 69 70 74)
//  input bit  62 used   3 times (syndrom bits 66 67 71)
//  input bit  63 used   3 times (syndrom bits 63 64 68)
//  input bit  64 used   3 times (syndrom bits 60 61 65)
//  input bit  65 used   3 times (syndrom bits 57 58 62)
//  input bit  66 used   3 times (syndrom bits 54 55 59)
//  input bit  67 used   3 times (syndrom bits 51 52 56)
//  input bit  68 used   3 times (syndrom bits 48 49 53)
//  input bit  69 used   3 times (syndrom bits 45 46 50)
//  input bit  70 used   3 times (syndrom bits 42 43 47)
//  input bit  71 used   3 times (syndrom bits 39 40 44)
//  input bit  72 used   3 times (syndrom bits 36 37 41)
//  input bit  73 used   3 times (syndrom bits 33 34 38)
//  input bit  74 used   3 times (syndrom bits 30 31 35)
//  input bit  75 used   3 times (syndrom bits 27 28 32)
//  input bit  76 used   3 times (syndrom bits 24 25 29)
//  input bit  77 used   3 times (syndrom bits 21 22 26)
//  input bit  78 used   3 times (syndrom bits 18 19 23)
//  input bit  79 used   3 times (syndrom bits 15 16 20)
//  input bit  80 used   3 times (syndrom bits 12 13 17)
//  input bit  81 used   3 times (syndrom bits 9 10 14)
//  input bit  82 used   3 times (syndrom bits 6 7 11)
//  input bit  83 used   3 times (syndrom bits 3 4 8)
//  input bit  84 used   3 times (syndrom bits 0 1 5)
//  input bit  85 used   3 times (syndrom bits 0 2 5)
//  input bit  86 used   3 times (syndrom bits 1 2 8)
//  input bit  87 used   3 times (syndrom bits 3 4 11)
//  input bit  88 used   3 times (syndrom bits 6 7 14)
//  input bit  89 used   3 times (syndrom bits 9 10 17)
//  input bit  90 used   3 times (syndrom bits 12 13 20)
//  input bit  91 used   3 times (syndrom bits 15 16 23)
//  input bit  92 used   3 times (syndrom bits 18 19 26)
//  input bit  93 used   3 times (syndrom bits 21 22 29)
//  input bit  94 used   3 times (syndrom bits 24 25 32)
//  input bit  95 used   3 times (syndrom bits 27 28 35)
//  input bit  96 used   3 times (syndrom bits 30 31 38)
//  input bit  97 used   3 times (syndrom bits 33 34 41)
//  input bit  98 used   3 times (syndrom bits 36 37 44)
//  input bit  99 used   3 times (syndrom bits 39 40 47)
//  input bit 100 used   3 times (syndrom bits 42 43 50)
//  input bit 101 used   3 times (syndrom bits 45 46 53)
//  input bit 102 used   3 times (syndrom bits 48 49 56)
//  input bit 103 used   3 times (syndrom bits 51 52 59)
//  input bit 104 used   3 times (syndrom bits 54 55 62)
//  input bit 105 used   3 times (syndrom bits 57 58 65)
//  input bit 106 used   3 times (syndrom bits 60 61 68)
//  input bit 107 used   3 times (syndrom bits 63 64 71)
//  input bit 108 used   3 times (syndrom bits 66 67 74)
//  input bit 109 used   3 times (syndrom bits 69 70 77)
//  input bit 110 used   3 times (syndrom bits 72 73 80)
//  input bit 111 used   3 times (syndrom bits 75 76 83)
//  input bit 112 used   3 times (syndrom bits 78 79 86)
//  input bit 113 used   3 times (syndrom bits 81 82 89)
//  input bit 114 used   3 times (syndrom bits 84 85 92)
//  input bit 115 used   3 times (syndrom bits 87 88 95)
//  input bit 116 used   3 times (syndrom bits 90 91 98)
//  input bit 117 used   3 times (syndrom bits 93 94 101)
//  input bit 118 used   3 times (syndrom bits 96 97 104)
//  input bit 119 used   3 times (syndrom bits 99 100 107)
//  input bit 120 used   3 times (syndrom bits 102 103 110)
//  input bit 121 used   3 times (syndrom bits 105 106 113)
//  input bit 122 used   3 times (syndrom bits 108 109 116)
//  input bit 123 used   3 times (syndrom bits 111 112 119)
//  input bit 124 used   3 times (syndrom bits 114 115 122)
//  input bit 125 used   3 times (syndrom bits 117 118 125)
//  input bit 126 used   3 times (syndrom bits 120 121 126)
//  input bit 127 used   3 times (syndrom bits 123 124 127)
function [128-1:0] extended_hamming_code_256_128_f;
    input [128-1:0] in;
    reg [128-1:0] syndrom;
    begin
        syndrom[  0] = in[  0]^in[ 84]^in[ 85];//3 inputs
        syndrom[  1] = in[  0]^in[ 84]^in[ 86];//3 inputs
        syndrom[  2] = in[  0]^in[ 85]^in[ 86];//3 inputs
        syndrom[  3] = in[  1]^in[ 83]^in[ 87];//3 inputs
        syndrom[  4] = in[  1]^in[ 83]^in[ 87];//3 inputs
        syndrom[  5] = in[  1]^in[ 84]^in[ 85];//3 inputs
        syndrom[  6] = in[  2]^in[ 82]^in[ 88];//3 inputs
        syndrom[  7] = in[  2]^in[ 82]^in[ 88];//3 inputs
        syndrom[  8] = in[  2]^in[ 83]^in[ 86];//3 inputs
        syndrom[  9] = in[  3]^in[ 81]^in[ 89];//3 inputs
        syndrom[ 10] = in[  3]^in[ 81]^in[ 89];//3 inputs
        syndrom[ 11] = in[  3]^in[ 82]^in[ 87];//3 inputs
        syndrom[ 12] = in[  4]^in[ 80]^in[ 90];//3 inputs
        syndrom[ 13] = in[  4]^in[ 80]^in[ 90];//3 inputs
        syndrom[ 14] = in[  4]^in[ 81]^in[ 88];//3 inputs
        syndrom[ 15] = in[  5]^in[ 79]^in[ 91];//3 inputs
        syndrom[ 16] = in[  5]^in[ 79]^in[ 91];//3 inputs
        syndrom[ 17] = in[  5]^in[ 80]^in[ 89];//3 inputs
        syndrom[ 18] = in[  6]^in[ 78]^in[ 92];//3 inputs
        syndrom[ 19] = in[  6]^in[ 78]^in[ 92];//3 inputs
        syndrom[ 20] = in[  6]^in[ 79]^in[ 90];//3 inputs
        syndrom[ 21] = in[  7]^in[ 77]^in[ 93];//3 inputs
        syndrom[ 22] = in[  7]^in[ 77]^in[ 93];//3 inputs
        syndrom[ 23] = in[  7]^in[ 78]^in[ 91];//3 inputs
        syndrom[ 24] = in[  8]^in[ 76]^in[ 94];//3 inputs
        syndrom[ 25] = in[  8]^in[ 76]^in[ 94];//3 inputs
        syndrom[ 26] = in[  8]^in[ 77]^in[ 92];//3 inputs
        syndrom[ 27] = in[  9]^in[ 75]^in[ 95];//3 inputs
        syndrom[ 28] = in[  9]^in[ 75]^in[ 95];//3 inputs
        syndrom[ 29] = in[  9]^in[ 76]^in[ 93];//3 inputs
        syndrom[ 30] = in[ 10]^in[ 74]^in[ 96];//3 inputs
        syndrom[ 31] = in[ 10]^in[ 74]^in[ 96];//3 inputs
        syndrom[ 32] = in[ 10]^in[ 75]^in[ 94];//3 inputs
        syndrom[ 33] = in[ 11]^in[ 73]^in[ 97];//3 inputs
        syndrom[ 34] = in[ 11]^in[ 73]^in[ 97];//3 inputs
        syndrom[ 35] = in[ 11]^in[ 74]^in[ 95];//3 inputs
        syndrom[ 36] = in[ 12]^in[ 72]^in[ 98];//3 inputs
        syndrom[ 37] = in[ 12]^in[ 72]^in[ 98];//3 inputs
        syndrom[ 38] = in[ 12]^in[ 73]^in[ 96];//3 inputs
        syndrom[ 39] = in[ 13]^in[ 71]^in[ 99];//3 inputs
        syndrom[ 40] = in[ 13]^in[ 71]^in[ 99];//3 inputs
        syndrom[ 41] = in[ 13]^in[ 72]^in[ 97];//3 inputs
        syndrom[ 42] = in[ 14]^in[ 70]^in[100];//3 inputs
        syndrom[ 43] = in[ 14]^in[ 70]^in[100];//3 inputs
        syndrom[ 44] = in[ 14]^in[ 71]^in[ 98];//3 inputs
        syndrom[ 45] = in[ 15]^in[ 69]^in[101];//3 inputs
        syndrom[ 46] = in[ 15]^in[ 69]^in[101];//3 inputs
        syndrom[ 47] = in[ 15]^in[ 70]^in[ 99];//3 inputs
        syndrom[ 48] = in[ 16]^in[ 68]^in[102];//3 inputs
        syndrom[ 49] = in[ 16]^in[ 68]^in[102];//3 inputs
        syndrom[ 50] = in[ 16]^in[ 69]^in[100];//3 inputs
        syndrom[ 51] = in[ 17]^in[ 67]^in[103];//3 inputs
        syndrom[ 52] = in[ 17]^in[ 67]^in[103];//3 inputs
        syndrom[ 53] = in[ 17]^in[ 68]^in[101];//3 inputs
        syndrom[ 54] = in[ 18]^in[ 66]^in[104];//3 inputs
        syndrom[ 55] = in[ 18]^in[ 66]^in[104];//3 inputs
        syndrom[ 56] = in[ 18]^in[ 67]^in[102];//3 inputs
        syndrom[ 57] = in[ 19]^in[ 65]^in[105];//3 inputs
        syndrom[ 58] = in[ 19]^in[ 65]^in[105];//3 inputs
        syndrom[ 59] = in[ 19]^in[ 66]^in[103];//3 inputs
        syndrom[ 60] = in[ 20]^in[ 64]^in[106];//3 inputs
        syndrom[ 61] = in[ 20]^in[ 64]^in[106];//3 inputs
        syndrom[ 62] = in[ 20]^in[ 65]^in[104];//3 inputs
        syndrom[ 63] = in[ 21]^in[ 63]^in[107];//3 inputs
        syndrom[ 64] = in[ 21]^in[ 63]^in[107];//3 inputs
        syndrom[ 65] = in[ 21]^in[ 64]^in[105];//3 inputs
        syndrom[ 66] = in[ 22]^in[ 62]^in[108];//3 inputs
        syndrom[ 67] = in[ 22]^in[ 62]^in[108];//3 inputs
        syndrom[ 68] = in[ 22]^in[ 63]^in[106];//3 inputs
        syndrom[ 69] = in[ 23]^in[ 61]^in[109];//3 inputs
        syndrom[ 70] = in[ 23]^in[ 61]^in[109];//3 inputs
        syndrom[ 71] = in[ 23]^in[ 62]^in[107];//3 inputs
        syndrom[ 72] = in[ 24]^in[ 60]^in[110];//3 inputs
        syndrom[ 73] = in[ 24]^in[ 60]^in[110];//3 inputs
        syndrom[ 74] = in[ 24]^in[ 61]^in[108];//3 inputs
        syndrom[ 75] = in[ 25]^in[ 59]^in[111];//3 inputs
        syndrom[ 76] = in[ 25]^in[ 59]^in[111];//3 inputs
        syndrom[ 77] = in[ 25]^in[ 60]^in[109];//3 inputs
        syndrom[ 78] = in[ 26]^in[ 58]^in[112];//3 inputs
        syndrom[ 79] = in[ 26]^in[ 58]^in[112];//3 inputs
        syndrom[ 80] = in[ 26]^in[ 59]^in[110];//3 inputs
        syndrom[ 81] = in[ 27]^in[ 57]^in[113];//3 inputs
        syndrom[ 82] = in[ 27]^in[ 57]^in[113];//3 inputs
        syndrom[ 83] = in[ 27]^in[ 58]^in[111];//3 inputs
        syndrom[ 84] = in[ 28]^in[ 56]^in[114];//3 inputs
        syndrom[ 85] = in[ 28]^in[ 56]^in[114];//3 inputs
        syndrom[ 86] = in[ 28]^in[ 57]^in[112];//3 inputs
        syndrom[ 87] = in[ 29]^in[ 55]^in[115];//3 inputs
        syndrom[ 88] = in[ 29]^in[ 55]^in[115];//3 inputs
        syndrom[ 89] = in[ 29]^in[ 56]^in[113];//3 inputs
        syndrom[ 90] = in[ 30]^in[ 54]^in[116];//3 inputs
        syndrom[ 91] = in[ 30]^in[ 54]^in[116];//3 inputs
        syndrom[ 92] = in[ 30]^in[ 55]^in[114];//3 inputs
        syndrom[ 93] = in[ 31]^in[ 53]^in[117];//3 inputs
        syndrom[ 94] = in[ 31]^in[ 53]^in[117];//3 inputs
        syndrom[ 95] = in[ 31]^in[ 54]^in[115];//3 inputs
        syndrom[ 96] = in[ 32]^in[ 52]^in[118];//3 inputs
        syndrom[ 97] = in[ 32]^in[ 52]^in[118];//3 inputs
        syndrom[ 98] = in[ 32]^in[ 53]^in[116];//3 inputs
        syndrom[ 99] = in[ 33]^in[ 51]^in[119];//3 inputs
        syndrom[100] = in[ 33]^in[ 51]^in[119];//3 inputs
        syndrom[101] = in[ 33]^in[ 52]^in[117];//3 inputs
        syndrom[102] = in[ 34]^in[ 50]^in[120];//3 inputs
        syndrom[103] = in[ 34]^in[ 50]^in[120];//3 inputs
        syndrom[104] = in[ 34]^in[ 51]^in[118];//3 inputs
        syndrom[105] = in[ 35]^in[ 49]^in[121];//3 inputs
        syndrom[106] = in[ 35]^in[ 49]^in[121];//3 inputs
        syndrom[107] = in[ 35]^in[ 50]^in[119];//3 inputs
        syndrom[108] = in[ 36]^in[ 48]^in[122];//3 inputs
        syndrom[109] = in[ 36]^in[ 48]^in[122];//3 inputs
        syndrom[110] = in[ 36]^in[ 49]^in[120];//3 inputs
        syndrom[111] = in[ 37]^in[ 47]^in[123];//3 inputs
        syndrom[112] = in[ 37]^in[ 47]^in[123];//3 inputs
        syndrom[113] = in[ 37]^in[ 48]^in[121];//3 inputs
        syndrom[114] = in[ 38]^in[ 46]^in[124];//3 inputs
        syndrom[115] = in[ 38]^in[ 46]^in[124];//3 inputs
        syndrom[116] = in[ 38]^in[ 47]^in[122];//3 inputs
        syndrom[117] = in[ 39]^in[ 45]^in[125];//3 inputs
        syndrom[118] = in[ 39]^in[ 45]^in[125];//3 inputs
        syndrom[119] = in[ 39]^in[ 46]^in[123];//3 inputs
        syndrom[120] = in[ 40]^in[ 44]^in[126];//3 inputs
        syndrom[121] = in[ 40]^in[ 44]^in[126];//3 inputs
        syndrom[122] = in[ 40]^in[ 45]^in[124];//3 inputs
        syndrom[123] = in[ 41]^in[ 42]^in[127];//3 inputs
        syndrom[124] = in[ 41]^in[ 43]^in[127];//3 inputs
        syndrom[125] = in[ 41]^in[ 44]^in[125];//3 inputs
        syndrom[126] = in[ 42]^in[ 43]^in[126];//3 inputs
        syndrom[127] = in[ 42]^in[ 43]^in[127];//3 inputs
        extended_hamming_code_256_128_f = syndrom;
    end
endfunction
wire [128-1:0] stored_data_edc = extended_hamming_code_256_128_f(i_stored_data);
wire [128-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_128_min_delay (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [128-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [128-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [128-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_256_128_f
//Compute 128 bits Error Detection Code from a 128 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used   3 times (syndrom bits 0 1 2)
//  input bit   1 used   3 times (syndrom bits 3 4 5)
//  input bit   2 used   3 times (syndrom bits 6 7 8)
//  input bit   3 used   3 times (syndrom bits 9 10 11)
//  input bit   4 used   3 times (syndrom bits 12 13 14)
//  input bit   5 used   3 times (syndrom bits 15 16 17)
//  input bit   6 used   3 times (syndrom bits 18 19 20)
//  input bit   7 used   3 times (syndrom bits 21 22 23)
//  input bit   8 used   3 times (syndrom bits 24 25 26)
//  input bit   9 used   3 times (syndrom bits 27 28 29)
//  input bit  10 used   3 times (syndrom bits 30 31 32)
//  input bit  11 used   3 times (syndrom bits 33 34 35)
//  input bit  12 used   3 times (syndrom bits 36 37 38)
//  input bit  13 used   3 times (syndrom bits 39 40 41)
//  input bit  14 used   3 times (syndrom bits 42 43 44)
//  input bit  15 used   3 times (syndrom bits 45 46 47)
//  input bit  16 used   3 times (syndrom bits 48 49 50)
//  input bit  17 used   3 times (syndrom bits 51 52 53)
//  input bit  18 used   3 times (syndrom bits 54 55 56)
//  input bit  19 used   3 times (syndrom bits 57 58 59)
//  input bit  20 used   3 times (syndrom bits 60 61 62)
//  input bit  21 used   3 times (syndrom bits 63 64 65)
//  input bit  22 used   3 times (syndrom bits 66 67 68)
//  input bit  23 used   3 times (syndrom bits 69 70 71)
//  input bit  24 used   3 times (syndrom bits 72 73 74)
//  input bit  25 used   3 times (syndrom bits 75 76 77)
//  input bit  26 used   3 times (syndrom bits 78 79 80)
//  input bit  27 used   3 times (syndrom bits 81 82 83)
//  input bit  28 used   3 times (syndrom bits 84 85 86)
//  input bit  29 used   3 times (syndrom bits 87 88 89)
//  input bit  30 used   3 times (syndrom bits 90 91 92)
//  input bit  31 used   3 times (syndrom bits 93 94 95)
//  input bit  32 used   3 times (syndrom bits 96 97 98)
//  input bit  33 used   3 times (syndrom bits 99 100 101)
//  input bit  34 used   3 times (syndrom bits 102 103 104)
//  input bit  35 used   3 times (syndrom bits 105 106 107)
//  input bit  36 used   3 times (syndrom bits 108 109 110)
//  input bit  37 used   3 times (syndrom bits 111 112 113)
//  input bit  38 used   3 times (syndrom bits 114 115 116)
//  input bit  39 used   3 times (syndrom bits 117 118 119)
//  input bit  40 used   3 times (syndrom bits 120 121 122)
//  input bit  41 used   3 times (syndrom bits 123 124 125)
//  input bit  42 used   3 times (syndrom bits 123 126 127)
//  input bit  43 used   3 times (syndrom bits 124 126 127)
//  input bit  44 used   3 times (syndrom bits 120 121 125)
//  input bit  45 used   3 times (syndrom bits 117 118 122)
//  input bit  46 used   3 times (syndrom bits 114 115 119)
//  input bit  47 used   3 times (syndrom bits 111 112 116)
//  input bit  48 used   3 times (syndrom bits 108 109 113)
//  input bit  49 used   3 times (syndrom bits 105 106 110)
//  input bit  50 used   3 times (syndrom bits 102 103 107)
//  input bit  51 used   3 times (syndrom bits 99 100 104)
//  input bit  52 used   3 times (syndrom bits 96 97 101)
//  input bit  53 used   3 times (syndrom bits 93 94 98)
//  input bit  54 used   3 times (syndrom bits 90 91 95)
//  input bit  55 used   3 times (syndrom bits 87 88 92)
//  input bit  56 used   3 times (syndrom bits 84 85 89)
//  input bit  57 used   3 times (syndrom bits 81 82 86)
//  input bit  58 used   3 times (syndrom bits 78 79 83)
//  input bit  59 used   3 times (syndrom bits 75 76 80)
//  input bit  60 used   3 times (syndrom bits 72 73 77)
//  input bit  61 used   3 times (syndrom bits 69 70 74)
//  input bit  62 used   3 times (syndrom bits 66 67 71)
//  input bit  63 used   3 times (syndrom bits 63 64 68)
//  input bit  64 used   3 times (syndrom bits 60 61 65)
//  input bit  65 used   3 times (syndrom bits 57 58 62)
//  input bit  66 used   3 times (syndrom bits 54 55 59)
//  input bit  67 used   3 times (syndrom bits 51 52 56)
//  input bit  68 used   3 times (syndrom bits 48 49 53)
//  input bit  69 used   3 times (syndrom bits 45 46 50)
//  input bit  70 used   3 times (syndrom bits 42 43 47)
//  input bit  71 used   3 times (syndrom bits 39 40 44)
//  input bit  72 used   3 times (syndrom bits 36 37 41)
//  input bit  73 used   3 times (syndrom bits 33 34 38)
//  input bit  74 used   3 times (syndrom bits 30 31 35)
//  input bit  75 used   3 times (syndrom bits 27 28 32)
//  input bit  76 used   3 times (syndrom bits 24 25 29)
//  input bit  77 used   3 times (syndrom bits 21 22 26)
//  input bit  78 used   3 times (syndrom bits 18 19 23)
//  input bit  79 used   3 times (syndrom bits 15 16 20)
//  input bit  80 used   3 times (syndrom bits 12 13 17)
//  input bit  81 used   3 times (syndrom bits 9 10 14)
//  input bit  82 used   3 times (syndrom bits 6 7 11)
//  input bit  83 used   3 times (syndrom bits 3 4 8)
//  input bit  84 used   3 times (syndrom bits 0 1 5)
//  input bit  85 used   3 times (syndrom bits 0 2 5)
//  input bit  86 used   3 times (syndrom bits 1 2 8)
//  input bit  87 used   3 times (syndrom bits 3 4 11)
//  input bit  88 used   3 times (syndrom bits 6 7 14)
//  input bit  89 used   3 times (syndrom bits 9 10 17)
//  input bit  90 used   3 times (syndrom bits 12 13 20)
//  input bit  91 used   3 times (syndrom bits 15 16 23)
//  input bit  92 used   3 times (syndrom bits 18 19 26)
//  input bit  93 used   3 times (syndrom bits 21 22 29)
//  input bit  94 used   3 times (syndrom bits 24 25 32)
//  input bit  95 used   3 times (syndrom bits 27 28 35)
//  input bit  96 used   3 times (syndrom bits 30 31 38)
//  input bit  97 used   3 times (syndrom bits 33 34 41)
//  input bit  98 used   3 times (syndrom bits 36 37 44)
//  input bit  99 used   3 times (syndrom bits 39 40 47)
//  input bit 100 used   3 times (syndrom bits 42 43 50)
//  input bit 101 used   3 times (syndrom bits 45 46 53)
//  input bit 102 used   3 times (syndrom bits 48 49 56)
//  input bit 103 used   3 times (syndrom bits 51 52 59)
//  input bit 104 used   3 times (syndrom bits 54 55 62)
//  input bit 105 used   3 times (syndrom bits 57 58 65)
//  input bit 106 used   3 times (syndrom bits 60 61 68)
//  input bit 107 used   3 times (syndrom bits 63 64 71)
//  input bit 108 used   3 times (syndrom bits 66 67 74)
//  input bit 109 used   3 times (syndrom bits 69 70 77)
//  input bit 110 used   3 times (syndrom bits 72 73 80)
//  input bit 111 used   3 times (syndrom bits 75 76 83)
//  input bit 112 used   3 times (syndrom bits 78 79 86)
//  input bit 113 used   3 times (syndrom bits 81 82 89)
//  input bit 114 used   3 times (syndrom bits 84 85 92)
//  input bit 115 used   3 times (syndrom bits 87 88 95)
//  input bit 116 used   3 times (syndrom bits 90 91 98)
//  input bit 117 used   3 times (syndrom bits 93 94 101)
//  input bit 118 used   3 times (syndrom bits 96 97 104)
//  input bit 119 used   3 times (syndrom bits 99 100 107)
//  input bit 120 used   3 times (syndrom bits 102 103 110)
//  input bit 121 used   3 times (syndrom bits 105 106 113)
//  input bit 122 used   3 times (syndrom bits 108 109 116)
//  input bit 123 used   3 times (syndrom bits 111 112 119)
//  input bit 124 used   3 times (syndrom bits 114 115 122)
//  input bit 125 used   3 times (syndrom bits 117 118 125)
//  input bit 126 used   3 times (syndrom bits 120 121 126)
//  input bit 127 used   3 times (syndrom bits 123 124 127)
function [128-1:0] extended_hamming_code_256_128_f;
    input [128-1:0] in;
    reg [128-1:0] syndrom;
    begin
        syndrom[  0] = in[  0]^in[ 84]^in[ 85];//3 inputs
        syndrom[  1] = in[  0]^in[ 84]^in[ 86];//3 inputs
        syndrom[  2] = in[  0]^in[ 85]^in[ 86];//3 inputs
        syndrom[  3] = in[  1]^in[ 83]^in[ 87];//3 inputs
        syndrom[  4] = in[  1]^in[ 83]^in[ 87];//3 inputs
        syndrom[  5] = in[  1]^in[ 84]^in[ 85];//3 inputs
        syndrom[  6] = in[  2]^in[ 82]^in[ 88];//3 inputs
        syndrom[  7] = in[  2]^in[ 82]^in[ 88];//3 inputs
        syndrom[  8] = in[  2]^in[ 83]^in[ 86];//3 inputs
        syndrom[  9] = in[  3]^in[ 81]^in[ 89];//3 inputs
        syndrom[ 10] = in[  3]^in[ 81]^in[ 89];//3 inputs
        syndrom[ 11] = in[  3]^in[ 82]^in[ 87];//3 inputs
        syndrom[ 12] = in[  4]^in[ 80]^in[ 90];//3 inputs
        syndrom[ 13] = in[  4]^in[ 80]^in[ 90];//3 inputs
        syndrom[ 14] = in[  4]^in[ 81]^in[ 88];//3 inputs
        syndrom[ 15] = in[  5]^in[ 79]^in[ 91];//3 inputs
        syndrom[ 16] = in[  5]^in[ 79]^in[ 91];//3 inputs
        syndrom[ 17] = in[  5]^in[ 80]^in[ 89];//3 inputs
        syndrom[ 18] = in[  6]^in[ 78]^in[ 92];//3 inputs
        syndrom[ 19] = in[  6]^in[ 78]^in[ 92];//3 inputs
        syndrom[ 20] = in[  6]^in[ 79]^in[ 90];//3 inputs
        syndrom[ 21] = in[  7]^in[ 77]^in[ 93];//3 inputs
        syndrom[ 22] = in[  7]^in[ 77]^in[ 93];//3 inputs
        syndrom[ 23] = in[  7]^in[ 78]^in[ 91];//3 inputs
        syndrom[ 24] = in[  8]^in[ 76]^in[ 94];//3 inputs
        syndrom[ 25] = in[  8]^in[ 76]^in[ 94];//3 inputs
        syndrom[ 26] = in[  8]^in[ 77]^in[ 92];//3 inputs
        syndrom[ 27] = in[  9]^in[ 75]^in[ 95];//3 inputs
        syndrom[ 28] = in[  9]^in[ 75]^in[ 95];//3 inputs
        syndrom[ 29] = in[  9]^in[ 76]^in[ 93];//3 inputs
        syndrom[ 30] = in[ 10]^in[ 74]^in[ 96];//3 inputs
        syndrom[ 31] = in[ 10]^in[ 74]^in[ 96];//3 inputs
        syndrom[ 32] = in[ 10]^in[ 75]^in[ 94];//3 inputs
        syndrom[ 33] = in[ 11]^in[ 73]^in[ 97];//3 inputs
        syndrom[ 34] = in[ 11]^in[ 73]^in[ 97];//3 inputs
        syndrom[ 35] = in[ 11]^in[ 74]^in[ 95];//3 inputs
        syndrom[ 36] = in[ 12]^in[ 72]^in[ 98];//3 inputs
        syndrom[ 37] = in[ 12]^in[ 72]^in[ 98];//3 inputs
        syndrom[ 38] = in[ 12]^in[ 73]^in[ 96];//3 inputs
        syndrom[ 39] = in[ 13]^in[ 71]^in[ 99];//3 inputs
        syndrom[ 40] = in[ 13]^in[ 71]^in[ 99];//3 inputs
        syndrom[ 41] = in[ 13]^in[ 72]^in[ 97];//3 inputs
        syndrom[ 42] = in[ 14]^in[ 70]^in[100];//3 inputs
        syndrom[ 43] = in[ 14]^in[ 70]^in[100];//3 inputs
        syndrom[ 44] = in[ 14]^in[ 71]^in[ 98];//3 inputs
        syndrom[ 45] = in[ 15]^in[ 69]^in[101];//3 inputs
        syndrom[ 46] = in[ 15]^in[ 69]^in[101];//3 inputs
        syndrom[ 47] = in[ 15]^in[ 70]^in[ 99];//3 inputs
        syndrom[ 48] = in[ 16]^in[ 68]^in[102];//3 inputs
        syndrom[ 49] = in[ 16]^in[ 68]^in[102];//3 inputs
        syndrom[ 50] = in[ 16]^in[ 69]^in[100];//3 inputs
        syndrom[ 51] = in[ 17]^in[ 67]^in[103];//3 inputs
        syndrom[ 52] = in[ 17]^in[ 67]^in[103];//3 inputs
        syndrom[ 53] = in[ 17]^in[ 68]^in[101];//3 inputs
        syndrom[ 54] = in[ 18]^in[ 66]^in[104];//3 inputs
        syndrom[ 55] = in[ 18]^in[ 66]^in[104];//3 inputs
        syndrom[ 56] = in[ 18]^in[ 67]^in[102];//3 inputs
        syndrom[ 57] = in[ 19]^in[ 65]^in[105];//3 inputs
        syndrom[ 58] = in[ 19]^in[ 65]^in[105];//3 inputs
        syndrom[ 59] = in[ 19]^in[ 66]^in[103];//3 inputs
        syndrom[ 60] = in[ 20]^in[ 64]^in[106];//3 inputs
        syndrom[ 61] = in[ 20]^in[ 64]^in[106];//3 inputs
        syndrom[ 62] = in[ 20]^in[ 65]^in[104];//3 inputs
        syndrom[ 63] = in[ 21]^in[ 63]^in[107];//3 inputs
        syndrom[ 64] = in[ 21]^in[ 63]^in[107];//3 inputs
        syndrom[ 65] = in[ 21]^in[ 64]^in[105];//3 inputs
        syndrom[ 66] = in[ 22]^in[ 62]^in[108];//3 inputs
        syndrom[ 67] = in[ 22]^in[ 62]^in[108];//3 inputs
        syndrom[ 68] = in[ 22]^in[ 63]^in[106];//3 inputs
        syndrom[ 69] = in[ 23]^in[ 61]^in[109];//3 inputs
        syndrom[ 70] = in[ 23]^in[ 61]^in[109];//3 inputs
        syndrom[ 71] = in[ 23]^in[ 62]^in[107];//3 inputs
        syndrom[ 72] = in[ 24]^in[ 60]^in[110];//3 inputs
        syndrom[ 73] = in[ 24]^in[ 60]^in[110];//3 inputs
        syndrom[ 74] = in[ 24]^in[ 61]^in[108];//3 inputs
        syndrom[ 75] = in[ 25]^in[ 59]^in[111];//3 inputs
        syndrom[ 76] = in[ 25]^in[ 59]^in[111];//3 inputs
        syndrom[ 77] = in[ 25]^in[ 60]^in[109];//3 inputs
        syndrom[ 78] = in[ 26]^in[ 58]^in[112];//3 inputs
        syndrom[ 79] = in[ 26]^in[ 58]^in[112];//3 inputs
        syndrom[ 80] = in[ 26]^in[ 59]^in[110];//3 inputs
        syndrom[ 81] = in[ 27]^in[ 57]^in[113];//3 inputs
        syndrom[ 82] = in[ 27]^in[ 57]^in[113];//3 inputs
        syndrom[ 83] = in[ 27]^in[ 58]^in[111];//3 inputs
        syndrom[ 84] = in[ 28]^in[ 56]^in[114];//3 inputs
        syndrom[ 85] = in[ 28]^in[ 56]^in[114];//3 inputs
        syndrom[ 86] = in[ 28]^in[ 57]^in[112];//3 inputs
        syndrom[ 87] = in[ 29]^in[ 55]^in[115];//3 inputs
        syndrom[ 88] = in[ 29]^in[ 55]^in[115];//3 inputs
        syndrom[ 89] = in[ 29]^in[ 56]^in[113];//3 inputs
        syndrom[ 90] = in[ 30]^in[ 54]^in[116];//3 inputs
        syndrom[ 91] = in[ 30]^in[ 54]^in[116];//3 inputs
        syndrom[ 92] = in[ 30]^in[ 55]^in[114];//3 inputs
        syndrom[ 93] = in[ 31]^in[ 53]^in[117];//3 inputs
        syndrom[ 94] = in[ 31]^in[ 53]^in[117];//3 inputs
        syndrom[ 95] = in[ 31]^in[ 54]^in[115];//3 inputs
        syndrom[ 96] = in[ 32]^in[ 52]^in[118];//3 inputs
        syndrom[ 97] = in[ 32]^in[ 52]^in[118];//3 inputs
        syndrom[ 98] = in[ 32]^in[ 53]^in[116];//3 inputs
        syndrom[ 99] = in[ 33]^in[ 51]^in[119];//3 inputs
        syndrom[100] = in[ 33]^in[ 51]^in[119];//3 inputs
        syndrom[101] = in[ 33]^in[ 52]^in[117];//3 inputs
        syndrom[102] = in[ 34]^in[ 50]^in[120];//3 inputs
        syndrom[103] = in[ 34]^in[ 50]^in[120];//3 inputs
        syndrom[104] = in[ 34]^in[ 51]^in[118];//3 inputs
        syndrom[105] = in[ 35]^in[ 49]^in[121];//3 inputs
        syndrom[106] = in[ 35]^in[ 49]^in[121];//3 inputs
        syndrom[107] = in[ 35]^in[ 50]^in[119];//3 inputs
        syndrom[108] = in[ 36]^in[ 48]^in[122];//3 inputs
        syndrom[109] = in[ 36]^in[ 48]^in[122];//3 inputs
        syndrom[110] = in[ 36]^in[ 49]^in[120];//3 inputs
        syndrom[111] = in[ 37]^in[ 47]^in[123];//3 inputs
        syndrom[112] = in[ 37]^in[ 47]^in[123];//3 inputs
        syndrom[113] = in[ 37]^in[ 48]^in[121];//3 inputs
        syndrom[114] = in[ 38]^in[ 46]^in[124];//3 inputs
        syndrom[115] = in[ 38]^in[ 46]^in[124];//3 inputs
        syndrom[116] = in[ 38]^in[ 47]^in[122];//3 inputs
        syndrom[117] = in[ 39]^in[ 45]^in[125];//3 inputs
        syndrom[118] = in[ 39]^in[ 45]^in[125];//3 inputs
        syndrom[119] = in[ 39]^in[ 46]^in[123];//3 inputs
        syndrom[120] = in[ 40]^in[ 44]^in[126];//3 inputs
        syndrom[121] = in[ 40]^in[ 44]^in[126];//3 inputs
        syndrom[122] = in[ 40]^in[ 45]^in[124];//3 inputs
        syndrom[123] = in[ 41]^in[ 42]^in[127];//3 inputs
        syndrom[124] = in[ 41]^in[ 43]^in[127];//3 inputs
        syndrom[125] = in[ 41]^in[ 44]^in[125];//3 inputs
        syndrom[126] = in[ 42]^in[ 43]^in[126];//3 inputs
        syndrom[127] = in[ 42]^in[ 43]^in[127];//3 inputs
        extended_hamming_code_256_128_f = syndrom;
    end
endfunction
function [2+128-1:0] extended_hamming_code_256_128_f_correction_pattern_f;
    input [128-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [128-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {128{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {128{1'b0}};
			end	
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111: begin
				correction_pattern = {128{1'b0}};correction_pattern[  0]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  1]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  2]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  3]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  4]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  5]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  6]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  7]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  8]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  9]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 10]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 11]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 12]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 13]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 14]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 15]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 16]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 17]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 18]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 19]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 20]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 21]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 22]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 23]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 24]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 25]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 26]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 27]=1'b1;
			end
			128'b00000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 28]=1'b1;
			end
			128'b00000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 29]=1'b1;
			end
			128'b00000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 30]=1'b1;
			end
			128'b00000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 31]=1'b1;
			end
			128'b00000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 32]=1'b1;
			end
			128'b00000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 33]=1'b1;
			end
			128'b00000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 34]=1'b1;
			end
			128'b00000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 35]=1'b1;
			end
			128'b00000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 36]=1'b1;
			end
			128'b00000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 37]=1'b1;
			end
			128'b00000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 38]=1'b1;
			end
			128'b00000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 39]=1'b1;
			end
			128'b00000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 40]=1'b1;
			end
			128'b00111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 41]=1'b1;
			end
			128'b11001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 42]=1'b1;
			end
			128'b11010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 43]=1'b1;
			end
			128'b00100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 44]=1'b1;
			end
			128'b00000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 45]=1'b1;
			end
			128'b00000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 46]=1'b1;
			end
			128'b00000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 47]=1'b1;
			end
			128'b00000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 48]=1'b1;
			end
			128'b00000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 49]=1'b1;
			end
			128'b00000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 50]=1'b1;
			end
			128'b00000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 51]=1'b1;
			end
			128'b00000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 52]=1'b1;
			end
			128'b00000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 53]=1'b1;
			end
			128'b00000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 54]=1'b1;
			end
			128'b00000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 55]=1'b1;
			end
			128'b00000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 56]=1'b1;
			end
			128'b00000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 57]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 58]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 59]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 60]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 61]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 62]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 63]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 64]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 65]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 66]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 67]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 68]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 69]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 70]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 71]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 72]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 73]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 74]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 75]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 76]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 77]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 78]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 79]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 80]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 81]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 82]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 83]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 84]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 85]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 86]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 87]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 88]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 89]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 90]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 91]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 92]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 93]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 94]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 95]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 96]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 97]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 98]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 99]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[100]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[101]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[102]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[103]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[104]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[105]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[106]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[107]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[108]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[109]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[110]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[111]=1'b1;
			end
			128'b00000000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[112]=1'b1;
			end
			128'b00000000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[113]=1'b1;
			end
			128'b00000000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[114]=1'b1;
			end
			128'b00000000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[115]=1'b1;
			end
			128'b00000000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[116]=1'b1;
			end
			128'b00000000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[117]=1'b1;
			end
			128'b00000000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[118]=1'b1;
			end
			128'b00000000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[119]=1'b1;
			end
			128'b00000000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[120]=1'b1;
			end
			128'b00000000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[121]=1'b1;
			end
			128'b00000000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[122]=1'b1;
			end
			128'b00000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[123]=1'b1;
			end
			128'b00000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[124]=1'b1;
			end
			128'b00100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[125]=1'b1;
			end
			128'b01000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[126]=1'b1;
			end
			128'b10011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[127]=1'b1;
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_256_128_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [128-1:0] stored_data_edc = extended_hamming_code_256_128_f(i_stored_data);
wire [128-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [128-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_256_128_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule


/////////////////////////////////////////////////////////////////////////////////////////////////
// *_balanced modules: balanced trade-off between logic depth and EDC width.
//EDC width is half of data's width or the minimum width + 1 for small input sizes.
/////////////////////////////////////////////////////////////////////////////////////////////////
module edc_hc_4_balanced (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: x x  (2 inputs)
//  syndrom[1]: x  x (2 inputs)
//  syndrom[2]:  xx  (2 inputs)
//  syndrom[3]:  x x (2 inputs)
//Input usage report:
//  input bit 0 used 2 times (syndrom bits 0 1)
//  input bit 1 used 2 times (syndrom bits 2 3)
//  input bit 2 used 2 times (syndrom bits 0 2)
//  input bit 3 used 2 times (syndrom bits 1 3)
function [4-1:0] hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[2];//2 inputs
        syndrom[1] = in[0]^in[3];//2 inputs
        syndrom[2] = in[1]^in[2];//2 inputs
        syndrom[3] = in[1]^in[3];//2 inputs
        hamming_code_8_4_f = syndrom;
    end
endfunction
wire [4-1:0] stored_data_edc = hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_4_balanced (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: xxx  (3 inputs)
//  syndrom[1]: xx x (3 inputs)
//  syndrom[2]: x xx (3 inputs)
//  syndrom[3]:  xxx (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 1 3)
//  input bit 2 used 3 times (syndrom bits 0 2 3)
//  input bit 3 used 3 times (syndrom bits 1 2 3)
function [4-1:0] extended_hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[2];//3 inputs
        syndrom[1] = in[0]^in[1]^in[3];//3 inputs
        syndrom[2] = in[0]^in[2]^in[3];//3 inputs
        syndrom[3] = in[1]^in[2]^in[3];//3 inputs
        extended_hamming_code_8_4_f = syndrom;
    end
endfunction
wire [4-1:0] stored_data_edc = extended_hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_4_balanced (
	input wire [4-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [4-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [4-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_8_4_f
//Compute 4 bits Error Detection Code from a 4 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16 valid code words out of 256 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[3]
//  syndrom[0]: xxx  (3 inputs)
//  syndrom[1]: xx x (3 inputs)
//  syndrom[2]: x xx (3 inputs)
//  syndrom[3]:  xxx (3 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 0 1 3)
//  input bit 2 used 3 times (syndrom bits 0 2 3)
//  input bit 3 used 3 times (syndrom bits 1 2 3)
function [4-1:0] extended_hamming_code_8_4_f;
    input [4-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[1]^in[2];//3 inputs
        syndrom[1] = in[0]^in[1]^in[3];//3 inputs
        syndrom[2] = in[0]^in[2]^in[3];//3 inputs
        syndrom[3] = in[1]^in[2]^in[3];//3 inputs
        extended_hamming_code_8_4_f = syndrom;
    end
endfunction
function [2+4-1:0] extended_hamming_code_8_4_f_correction_pattern_f;
    input [4-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [4-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {4{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			4'b0000: begin
				correctable_error = 1'b0;
				correction_pattern = {4{1'b0}};
			end	
			4'b0111: begin
				correction_pattern = {4{1'b0}};correction_pattern[0]=1'b1;
			end
			4'b1011: begin
				correction_pattern = {4{1'b0}};correction_pattern[1]=1'b1;
			end
			4'b1101: begin
				correction_pattern = {4{1'b0}};correction_pattern[2]=1'b1;
			end
			4'b1110: begin
				correction_pattern = {4{1'b0}};correction_pattern[3]=1'b1;
			end
			4'b0001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b0010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b0100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			4'b1000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {4{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_8_4_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [4-1:0] stored_data_edc = extended_hamming_code_8_4_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [4-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_8_4_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_8_balanced (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [4-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [4-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_12_8_f
//Compute 4 bits Error Detection Code from a 8 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 256 valid code words out of 4096 therefore 93% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: x x x  x (4 inputs)
//  syndrom[1]: x  x xxx (5 inputs)
//  syndrom[2]:  xx  xxx (5 inputs)
//  syndrom[3]:  x xx x  (4 inputs)
//Input usage report:
//  input bit 0 used 2 times (syndrom bits 0 1)
//  input bit 1 used 2 times (syndrom bits 2 3)
//  input bit 2 used 2 times (syndrom bits 0 2)
//  input bit 3 used 2 times (syndrom bits 1 3)
//  input bit 4 used 2 times (syndrom bits 0 3)
//  input bit 5 used 2 times (syndrom bits 1 2)
//  input bit 6 used 3 times (syndrom bits 1 2 3)
//  input bit 7 used 3 times (syndrom bits 0 1 2)
function [4-1:0] hamming_code_12_8_f;
    input [8-1:0] in;
    reg [4-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[2]^in[4]^in[7];//4 inputs
        syndrom[1] = in[0]^in[3]^in[5]^in[6]^in[7];//5 inputs
        syndrom[2] = in[1]^in[2]^in[5]^in[6]^in[7];//5 inputs
        syndrom[3] = in[1]^in[3]^in[4]^in[6];//4 inputs
        hamming_code_12_8_f = syndrom;
    end
endfunction
wire [4-1:0] stored_data_edc = hamming_code_12_8_f(i_stored_data);
wire [4-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_8_balanced (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_14_8_f
//Compute 6 bits Error Detection Code from a 8 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 256 valid code words out of 16384 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: x x  x x (4 inputs)
//  syndrom[1]: x  xx  x (4 inputs)
//  syndrom[2]: x  x xx  (4 inputs)
//  syndrom[3]:  xx x  x (4 inputs)
//  syndrom[4]:  xx  xx  (4 inputs)
//  syndrom[5]:  x xx x  (4 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 3 4 5)
//  input bit 2 used 3 times (syndrom bits 0 3 4)
//  input bit 3 used 3 times (syndrom bits 1 2 5)
//  input bit 4 used 3 times (syndrom bits 1 3 5)
//  input bit 5 used 3 times (syndrom bits 0 2 4)
//  input bit 6 used 3 times (syndrom bits 2 4 5)
//  input bit 7 used 3 times (syndrom bits 0 1 3)
function [6-1:0] extended_hamming_code_14_8_f;
    input [8-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[2]^in[5]^in[7];//4 inputs
        syndrom[1] = in[0]^in[3]^in[4]^in[7];//4 inputs
        syndrom[2] = in[0]^in[3]^in[5]^in[6];//4 inputs
        syndrom[3] = in[1]^in[2]^in[4]^in[7];//4 inputs
        syndrom[4] = in[1]^in[2]^in[5]^in[6];//4 inputs
        syndrom[5] = in[1]^in[3]^in[4]^in[6];//4 inputs
        extended_hamming_code_14_8_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = extended_hamming_code_14_8_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_8_balanced (
	input wire [8-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [8-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [8-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_14_8_f
//Compute 6 bits Error Detection Code from a 8 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 256 valid code words out of 16384 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[7]
//  syndrom[0]: x x  x x (4 inputs)
//  syndrom[1]: x  xx  x (4 inputs)
//  syndrom[2]: x  x xx  (4 inputs)
//  syndrom[3]:  xx x  x (4 inputs)
//  syndrom[4]:  xx  xx  (4 inputs)
//  syndrom[5]:  x xx x  (4 inputs)
//Input usage report:
//  input bit 0 used 3 times (syndrom bits 0 1 2)
//  input bit 1 used 3 times (syndrom bits 3 4 5)
//  input bit 2 used 3 times (syndrom bits 0 3 4)
//  input bit 3 used 3 times (syndrom bits 1 2 5)
//  input bit 4 used 3 times (syndrom bits 1 3 5)
//  input bit 5 used 3 times (syndrom bits 0 2 4)
//  input bit 6 used 3 times (syndrom bits 2 4 5)
//  input bit 7 used 3 times (syndrom bits 0 1 3)
function [6-1:0] extended_hamming_code_14_8_f;
    input [8-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[0]^in[2]^in[5]^in[7];//4 inputs
        syndrom[1] = in[0]^in[3]^in[4]^in[7];//4 inputs
        syndrom[2] = in[0]^in[3]^in[5]^in[6];//4 inputs
        syndrom[3] = in[1]^in[2]^in[4]^in[7];//4 inputs
        syndrom[4] = in[1]^in[2]^in[5]^in[6];//4 inputs
        syndrom[5] = in[1]^in[3]^in[4]^in[6];//4 inputs
        extended_hamming_code_14_8_f = syndrom;
    end
endfunction
function [2+8-1:0] extended_hamming_code_14_8_f_correction_pattern_f;
    input [6-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [8-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {8{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			6'b000000: begin
				correctable_error = 1'b0;
				correction_pattern = {8{1'b0}};
			end	
			6'b000111: begin
				correction_pattern = {8{1'b0}};correction_pattern[0]=1'b1;
			end
			6'b111000: begin
				correction_pattern = {8{1'b0}};correction_pattern[1]=1'b1;
			end
			6'b011001: begin
				correction_pattern = {8{1'b0}};correction_pattern[2]=1'b1;
			end
			6'b100110: begin
				correction_pattern = {8{1'b0}};correction_pattern[3]=1'b1;
			end
			6'b101010: begin
				correction_pattern = {8{1'b0}};correction_pattern[4]=1'b1;
			end
			6'b010101: begin
				correction_pattern = {8{1'b0}};correction_pattern[5]=1'b1;
			end
			6'b110100: begin
				correction_pattern = {8{1'b0}};correction_pattern[6]=1'b1;
			end
			6'b001011: begin
				correction_pattern = {8{1'b0}};correction_pattern[7]=1'b1;
			end
			6'b000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {8{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_14_8_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [6-1:0] stored_data_edc = extended_hamming_code_14_8_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [8-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_14_8_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_12_balanced (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_18_12_f
//Compute 6 bits Error Detection Code from a 12 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 262144 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[0]:      x  xx x (4 inputs)
//  syndrom[1]: x     xx  x  (4 inputs)
//  syndrom[2]:  x x    x x  (4 inputs)
//  syndrom[3]:  x  x x    x (4 inputs)
//  syndrom[4]:   xx   x x   (4 inputs)
//  syndrom[5]: x x xx       (4 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 1 5)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 2 4)
//  input bit  4 used 2 times (syndrom bits 3 5)
//  input bit  5 used 2 times (syndrom bits 0 5)
//  input bit  6 used 2 times (syndrom bits 1 3)
//  input bit  7 used 2 times (syndrom bits 1 4)
//  input bit  8 used 2 times (syndrom bits 0 2)
//  input bit  9 used 2 times (syndrom bits 0 4)
//  input bit 10 used 2 times (syndrom bits 1 2)
//  input bit 11 used 2 times (syndrom bits 0 3)
function [6-1:0] hamming_code_18_12_f;
    input [12-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 5]^in[ 8]^in[ 9]^in[11];//4 inputs
        syndrom[1] = in[ 0]^in[ 6]^in[ 7]^in[10];//4 inputs
        syndrom[2] = in[ 1]^in[ 3]^in[ 8]^in[10];//4 inputs
        syndrom[3] = in[ 1]^in[ 4]^in[ 6]^in[11];//4 inputs
        syndrom[4] = in[ 2]^in[ 3]^in[ 7]^in[ 9];//4 inputs
        syndrom[5] = in[ 0]^in[ 2]^in[ 4]^in[ 5];//4 inputs
        hamming_code_18_12_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = hamming_code_18_12_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_12_balanced (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_18_12_f
//Compute 6 bits Error Detection Code from a 12 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 262144 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[0]: x x  x xx x  (6 inputs)
//  syndrom[1]: x  xx  xx  x (6 inputs)
//  syndrom[2]: x  x xx  xx  (6 inputs)
//  syndrom[3]:  xx x  x xx  (6 inputs)
//  syndrom[4]:  xx  xx x  x (6 inputs)
//  syndrom[5]:  x xx x  x x (6 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
function [6-1:0] extended_hamming_code_18_12_f;
    input [12-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10];//6 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11];//6 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10];//6 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10];//6 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11];//6 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11];//6 inputs
        extended_hamming_code_18_12_f = syndrom;
    end
endfunction
wire [6-1:0] stored_data_edc = extended_hamming_code_18_12_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_12_balanced (
	input wire [12-1:0] i_write_data, // Data to write to storage
	output reg [6-1:0] o_write_edc, // EDC bits to write to storage
	input wire [12-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [6-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [12-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_18_12_f
//Compute 6 bits Error Detection Code from a 12 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4096 valid code words out of 262144 therefore 98% of errors are detected. 
//Dot graphic view: in[0]...in[11]
//  syndrom[0]: x x  x xx x  (6 inputs)
//  syndrom[1]: x  xx  xx  x (6 inputs)
//  syndrom[2]: x  x xx  xx  (6 inputs)
//  syndrom[3]:  xx x  x xx  (6 inputs)
//  syndrom[4]:  xx  xx x  x (6 inputs)
//  syndrom[5]:  x xx x  x x (6 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 0 3 4)
//  input bit  3 used 3 times (syndrom bits 1 2 5)
//  input bit  4 used 3 times (syndrom bits 1 3 5)
//  input bit  5 used 3 times (syndrom bits 0 2 4)
//  input bit  6 used 3 times (syndrom bits 2 4 5)
//  input bit  7 used 3 times (syndrom bits 0 1 3)
//  input bit  8 used 3 times (syndrom bits 0 1 4)
//  input bit  9 used 3 times (syndrom bits 2 3 5)
//  input bit 10 used 3 times (syndrom bits 0 2 3)
//  input bit 11 used 3 times (syndrom bits 1 4 5)
function [6-1:0] extended_hamming_code_18_12_f;
    input [12-1:0] in;
    reg [6-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 2]^in[ 5]^in[ 7]^in[ 8]^in[10];//6 inputs
        syndrom[1] = in[ 0]^in[ 3]^in[ 4]^in[ 7]^in[ 8]^in[11];//6 inputs
        syndrom[2] = in[ 0]^in[ 3]^in[ 5]^in[ 6]^in[ 9]^in[10];//6 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 4]^in[ 7]^in[ 9]^in[10];//6 inputs
        syndrom[4] = in[ 1]^in[ 2]^in[ 5]^in[ 6]^in[ 8]^in[11];//6 inputs
        syndrom[5] = in[ 1]^in[ 3]^in[ 4]^in[ 6]^in[ 9]^in[11];//6 inputs
        extended_hamming_code_18_12_f = syndrom;
    end
endfunction
function [2+12-1:0] extended_hamming_code_18_12_f_correction_pattern_f;
    input [6-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [12-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {12{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			6'b000000: begin
				correctable_error = 1'b0;
				correction_pattern = {12{1'b0}};
			end	
			6'b000111: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 0]=1'b1;
			end
			6'b111000: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 1]=1'b1;
			end
			6'b011001: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 2]=1'b1;
			end
			6'b100110: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 3]=1'b1;
			end
			6'b101010: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 4]=1'b1;
			end
			6'b010101: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 5]=1'b1;
			end
			6'b110100: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 6]=1'b1;
			end
			6'b001011: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 7]=1'b1;
			end
			6'b010011: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 8]=1'b1;
			end
			6'b101100: begin
				correction_pattern = {12{1'b0}};correction_pattern[ 9]=1'b1;
			end
			6'b001101: begin
				correction_pattern = {12{1'b0}};correction_pattern[10]=1'b1;
			end
			6'b110010: begin
				correction_pattern = {12{1'b0}};correction_pattern[11]=1'b1;
			end
			6'b000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			6'b100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {12{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_18_12_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [6-1:0] stored_data_edc = extended_hamming_code_18_12_f(i_stored_data);
wire [6-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [12-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_18_12_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_16_balanced (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_24_16_f
//Compute 8 bits Error Detection Code from a 16 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 16777216 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[0]: x     x x      x (4 inputs)
//  syndrom[1]: x      x x  x    (4 inputs)
//  syndrom[2]:  x    x  x   x   (4 inputs)
//  syndrom[3]:  x     xx     x  (4 inputs)
//  syndrom[4]:   x x     x    x (4 inputs)
//  syndrom[5]:   x  x     xx    (4 inputs)
//  syndrom[6]:    xx      x x   (4 inputs)
//  syndrom[7]:    x x    x   x  (4 inputs)
//Input usage report:
//  input bit  0 used 2 times (syndrom bits 0 1)
//  input bit  1 used 2 times (syndrom bits 2 3)
//  input bit  2 used 2 times (syndrom bits 4 5)
//  input bit  3 used 2 times (syndrom bits 6 7)
//  input bit  4 used 2 times (syndrom bits 4 6)
//  input bit  5 used 2 times (syndrom bits 5 7)
//  input bit  6 used 2 times (syndrom bits 0 2)
//  input bit  7 used 2 times (syndrom bits 1 3)
//  input bit  8 used 2 times (syndrom bits 0 3)
//  input bit  9 used 2 times (syndrom bits 1 2)
//  input bit 10 used 2 times (syndrom bits 4 7)
//  input bit 11 used 2 times (syndrom bits 5 6)
//  input bit 12 used 2 times (syndrom bits 1 5)
//  input bit 13 used 2 times (syndrom bits 2 6)
//  input bit 14 used 2 times (syndrom bits 3 7)
//  input bit 15 used 2 times (syndrom bits 0 4)
function [8-1:0] hamming_code_24_16_f;
    input [16-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 6]^in[ 8]^in[15];//4 inputs
        syndrom[1] = in[ 0]^in[ 7]^in[ 9]^in[12];//4 inputs
        syndrom[2] = in[ 1]^in[ 6]^in[ 9]^in[13];//4 inputs
        syndrom[3] = in[ 1]^in[ 7]^in[ 8]^in[14];//4 inputs
        syndrom[4] = in[ 2]^in[ 4]^in[10]^in[15];//4 inputs
        syndrom[5] = in[ 2]^in[ 5]^in[11]^in[12];//4 inputs
        syndrom[6] = in[ 3]^in[ 4]^in[11]^in[13];//4 inputs
        syndrom[7] = in[ 3]^in[ 5]^in[10]^in[14];//4 inputs
        hamming_code_24_16_f = syndrom;
    end
endfunction
wire [8-1:0] stored_data_edc = hamming_code_24_16_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_16_balanced (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_24_16_f
//Compute 8 bits Error Detection Code from a 16 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 16777216 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[0]: x   xx    xx   x (6 inputs)
//  syndrom[1]: x   x x  x  xx   (6 inputs)
//  syndrom[2]: x    xx x    xx  (6 inputs)
//  syndrom[3]:  xx    x xx    x (6 inputs)
//  syndrom[4]:  x x   xx   x x  (6 inputs)
//  syndrom[5]:  x  xx    xx  x  (6 inputs)
//  syndrom[6]:   xx  x  x x   x (6 inputs)
//  syndrom[7]:   xx   xx   xx   (6 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 6 7)
//  input bit  3 used 3 times (syndrom bits 4 6 7)
//  input bit  4 used 3 times (syndrom bits 0 1 5)
//  input bit  5 used 3 times (syndrom bits 0 2 5)
//  input bit  6 used 3 times (syndrom bits 1 2 6)
//  input bit  7 used 3 times (syndrom bits 3 4 7)
//  input bit  8 used 3 times (syndrom bits 2 4 7)
//  input bit  9 used 3 times (syndrom bits 1 3 6)
//  input bit 10 used 3 times (syndrom bits 0 3 5)
//  input bit 11 used 3 times (syndrom bits 0 5 6)
//  input bit 12 used 3 times (syndrom bits 1 4 7)
//  input bit 13 used 3 times (syndrom bits 1 2 7)
//  input bit 14 used 3 times (syndrom bits 2 4 5)
//  input bit 15 used 3 times (syndrom bits 0 3 6)
function [8-1:0] extended_hamming_code_24_16_f;
    input [16-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 5]^in[10]^in[11]^in[15];//6 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 6]^in[ 9]^in[12]^in[13];//6 inputs
        syndrom[2] = in[ 0]^in[ 5]^in[ 6]^in[ 8]^in[13]^in[14];//6 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 7]^in[ 9]^in[10]^in[15];//6 inputs
        syndrom[4] = in[ 1]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[14];//6 inputs
        syndrom[5] = in[ 1]^in[ 4]^in[ 5]^in[10]^in[11]^in[14];//6 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 6]^in[ 9]^in[11]^in[15];//6 inputs
        syndrom[7] = in[ 2]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[13];//6 inputs
        extended_hamming_code_24_16_f = syndrom;
    end
endfunction
wire [8-1:0] stored_data_edc = extended_hamming_code_24_16_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_16_balanced (
	input wire [16-1:0] i_write_data, // Data to write to storage
	output reg [8-1:0] o_write_edc, // EDC bits to write to storage
	input wire [16-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [8-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [16-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_24_16_f
//Compute 8 bits Error Detection Code from a 16 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 65536 valid code words out of 16777216 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[15]
//  syndrom[0]: x   xx    xx   x (6 inputs)
//  syndrom[1]: x   x x  x  xx   (6 inputs)
//  syndrom[2]: x    xx x    xx  (6 inputs)
//  syndrom[3]:  xx    x xx    x (6 inputs)
//  syndrom[4]:  x x   xx   x x  (6 inputs)
//  syndrom[5]:  x  xx    xx  x  (6 inputs)
//  syndrom[6]:   xx  x  x x   x (6 inputs)
//  syndrom[7]:   xx   xx   xx   (6 inputs)
//Input usage report:
//  input bit  0 used 3 times (syndrom bits 0 1 2)
//  input bit  1 used 3 times (syndrom bits 3 4 5)
//  input bit  2 used 3 times (syndrom bits 3 6 7)
//  input bit  3 used 3 times (syndrom bits 4 6 7)
//  input bit  4 used 3 times (syndrom bits 0 1 5)
//  input bit  5 used 3 times (syndrom bits 0 2 5)
//  input bit  6 used 3 times (syndrom bits 1 2 6)
//  input bit  7 used 3 times (syndrom bits 3 4 7)
//  input bit  8 used 3 times (syndrom bits 2 4 7)
//  input bit  9 used 3 times (syndrom bits 1 3 6)
//  input bit 10 used 3 times (syndrom bits 0 3 5)
//  input bit 11 used 3 times (syndrom bits 0 5 6)
//  input bit 12 used 3 times (syndrom bits 1 4 7)
//  input bit 13 used 3 times (syndrom bits 1 2 7)
//  input bit 14 used 3 times (syndrom bits 2 4 5)
//  input bit 15 used 3 times (syndrom bits 0 3 6)
function [8-1:0] extended_hamming_code_24_16_f;
    input [16-1:0] in;
    reg [8-1:0] syndrom;
    begin
        syndrom[0] = in[ 0]^in[ 4]^in[ 5]^in[10]^in[11]^in[15];//6 inputs
        syndrom[1] = in[ 0]^in[ 4]^in[ 6]^in[ 9]^in[12]^in[13];//6 inputs
        syndrom[2] = in[ 0]^in[ 5]^in[ 6]^in[ 8]^in[13]^in[14];//6 inputs
        syndrom[3] = in[ 1]^in[ 2]^in[ 7]^in[ 9]^in[10]^in[15];//6 inputs
        syndrom[4] = in[ 1]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[14];//6 inputs
        syndrom[5] = in[ 1]^in[ 4]^in[ 5]^in[10]^in[11]^in[14];//6 inputs
        syndrom[6] = in[ 2]^in[ 3]^in[ 6]^in[ 9]^in[11]^in[15];//6 inputs
        syndrom[7] = in[ 2]^in[ 3]^in[ 7]^in[ 8]^in[12]^in[13];//6 inputs
        extended_hamming_code_24_16_f = syndrom;
    end
endfunction
function [2+16-1:0] extended_hamming_code_24_16_f_correction_pattern_f;
    input [8-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [16-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {16{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			8'b00000000: begin
				correctable_error = 1'b0;
				correction_pattern = {16{1'b0}};
			end	
			8'b00000111: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 0]=1'b1;
			end
			8'b00111000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 1]=1'b1;
			end
			8'b11001000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 2]=1'b1;
			end
			8'b11010000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 3]=1'b1;
			end
			8'b00100011: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 4]=1'b1;
			end
			8'b00100101: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 5]=1'b1;
			end
			8'b01000110: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 6]=1'b1;
			end
			8'b10011000: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 7]=1'b1;
			end
			8'b10010100: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 8]=1'b1;
			end
			8'b01001010: begin
				correction_pattern = {16{1'b0}};correction_pattern[ 9]=1'b1;
			end
			8'b00101001: begin
				correction_pattern = {16{1'b0}};correction_pattern[10]=1'b1;
			end
			8'b01100001: begin
				correction_pattern = {16{1'b0}};correction_pattern[11]=1'b1;
			end
			8'b10010010: begin
				correction_pattern = {16{1'b0}};correction_pattern[12]=1'b1;
			end
			8'b10000110: begin
				correction_pattern = {16{1'b0}};correction_pattern[13]=1'b1;
			end
			8'b00110100: begin
				correction_pattern = {16{1'b0}};correction_pattern[14]=1'b1;
			end
			8'b01001001: begin
				correction_pattern = {16{1'b0}};correction_pattern[15]=1'b1;
			end
			8'b00000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b00100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b01000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			8'b10000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {16{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_24_16_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [8-1:0] stored_data_edc = extended_hamming_code_24_16_f(i_stored_data);
wire [8-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [16-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_24_16_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_20_balanced (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [10-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [10-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_30_20_f
//Compute 10 bits Error Detection Code from a 20 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 1073741824 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[ 0]: x        x  x  x     (4 inputs)
//  syndrom[ 1]: x         xx     x   (4 inputs)
//  syndrom[ 2]:  x     x    x   x    (4 inputs)
//  syndrom[ 3]:  x      x x        x (4 inputs)
//  syndrom[ 4]:   x    x   x      x  (4 inputs)
//  syndrom[ 5]:   xx    xx           (4 inputs)
//  syndrom[ 6]:      x       x    xx (4 inputs)
//  syndrom[ 7]:    x  x       xx     (4 inputs)
//  syndrom[ 8]:     xx        x x    (4 inputs)
//  syndrom[ 9]:     x x      x   x   (4 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 5 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 6 8)
//  input bit  6 used  2 times (syndrom bits 7 9)
//  input bit  7 used  2 times (syndrom bits 2 4)
//  input bit  8 used  2 times (syndrom bits 3 5)
//  input bit  9 used  2 times (syndrom bits 0 5)
//  input bit 10 used  2 times (syndrom bits 1 3)
//  input bit 11 used  2 times (syndrom bits 1 4)
//  input bit 12 used  2 times (syndrom bits 0 2)
//  input bit 13 used  2 times (syndrom bits 6 9)
//  input bit 14 used  2 times (syndrom bits 7 8)
//  input bit 15 used  2 times (syndrom bits 0 7)
//  input bit 16 used  2 times (syndrom bits 2 8)
//  input bit 17 used  2 times (syndrom bits 1 9)
//  input bit 18 used  2 times (syndrom bits 4 6)
//  input bit 19 used  2 times (syndrom bits 3 6)
function [10-1:0] hamming_code_30_20_f;
    input [20-1:0] in;
    reg [10-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 9]^in[12]^in[15];//4 inputs
        syndrom[ 1] = in[ 0]^in[10]^in[11]^in[17];//4 inputs
        syndrom[ 2] = in[ 1]^in[ 7]^in[12]^in[16];//4 inputs
        syndrom[ 3] = in[ 1]^in[ 8]^in[10]^in[19];//4 inputs
        syndrom[ 4] = in[ 2]^in[ 7]^in[11]^in[18];//4 inputs
        syndrom[ 5] = in[ 2]^in[ 3]^in[ 8]^in[ 9];//4 inputs
        syndrom[ 6] = in[ 5]^in[13]^in[18]^in[19];//4 inputs
        syndrom[ 7] = in[ 3]^in[ 6]^in[14]^in[15];//4 inputs
        syndrom[ 8] = in[ 4]^in[ 5]^in[14]^in[16];//4 inputs
        syndrom[ 9] = in[ 4]^in[ 6]^in[13]^in[17];//4 inputs
        hamming_code_30_20_f = syndrom;
    end
endfunction
wire [10-1:0] stored_data_edc = hamming_code_30_20_f(i_stored_data);
wire [10-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_20_balanced (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [10-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [10-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_30_20_f
//Compute 10 bits Error Detection Code from a 20 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 1073741824 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[ 0]: x    x  x x     xx   (6 inputs)
//  syndrom[ 1]: x     xx    xx     x (6 inputs)
//  syndrom[ 2]: x     xx    x x    x (6 inputs)
//  syndrom[ 3]:  x  x    xx     xx   (6 inputs)
//  syndrom[ 4]:  x   xx      xx   x  (6 inputs)
//  syndrom[ 5]:  x   x x     xx   x  (6 inputs)
//  syndrom[ 6]:   xx     x     x  xx (6 inputs)
//  syndrom[ 7]:   xx     xxxx        (6 inputs)
//  syndrom[ 8]:   x x   x  x   x x   (6 inputs)
//  syndrom[ 9]:    xx   x  x   xx    (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 6 7 9)
//  input bit  4 used  3 times (syndrom bits 3 8 9)
//  input bit  5 used  3 times (syndrom bits 0 4 5)
//  input bit  6 used  3 times (syndrom bits 1 2 4)
//  input bit  7 used  3 times (syndrom bits 1 2 5)
//  input bit  8 used  3 times (syndrom bits 0 8 9)
//  input bit  9 used  3 times (syndrom bits 3 6 7)
//  input bit 10 used  3 times (syndrom bits 0 3 7)
//  input bit 11 used  3 times (syndrom bits 7 8 9)
//  input bit 12 used  3 times (syndrom bits 1 2 7)
//  input bit 13 used  3 times (syndrom bits 1 4 5)
//  input bit 14 used  3 times (syndrom bits 2 4 5)
//  input bit 15 used  3 times (syndrom bits 6 8 9)
//  input bit 16 used  3 times (syndrom bits 0 3 9)
//  input bit 17 used  3 times (syndrom bits 0 3 8)
//  input bit 18 used  3 times (syndrom bits 4 5 6)
//  input bit 19 used  3 times (syndrom bits 1 2 6)
function [10-1:0] extended_hamming_code_30_20_f;
    input [20-1:0] in;
    reg [10-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 5]^in[ 8]^in[10]^in[16]^in[17];//6 inputs
        syndrom[ 1] = in[ 0]^in[ 6]^in[ 7]^in[12]^in[13]^in[19];//6 inputs
        syndrom[ 2] = in[ 0]^in[ 6]^in[ 7]^in[12]^in[14]^in[19];//6 inputs
        syndrom[ 3] = in[ 1]^in[ 4]^in[ 9]^in[10]^in[16]^in[17];//6 inputs
        syndrom[ 4] = in[ 1]^in[ 5]^in[ 6]^in[13]^in[14]^in[18];//6 inputs
        syndrom[ 5] = in[ 1]^in[ 5]^in[ 7]^in[13]^in[14]^in[18];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 3]^in[ 9]^in[15]^in[18]^in[19];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 3]^in[ 9]^in[10]^in[11]^in[12];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 4]^in[ 8]^in[11]^in[15]^in[17];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 4]^in[ 8]^in[11]^in[15]^in[16];//6 inputs
        extended_hamming_code_30_20_f = syndrom;
    end
endfunction
wire [10-1:0] stored_data_edc = extended_hamming_code_30_20_f(i_stored_data);
wire [10-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_20_balanced (
	input wire [20-1:0] i_write_data, // Data to write to storage
	output reg [10-1:0] o_write_edc, // EDC bits to write to storage
	input wire [20-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [10-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [20-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_30_20_f
//Compute 10 bits Error Detection Code from a 20 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1048576 valid code words out of 1073741824 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[19]
//  syndrom[ 0]: x    x  x x     xx   (6 inputs)
//  syndrom[ 1]: x     xx    xx     x (6 inputs)
//  syndrom[ 2]: x     xx    x x    x (6 inputs)
//  syndrom[ 3]:  x  x    xx     xx   (6 inputs)
//  syndrom[ 4]:  x   xx      xx   x  (6 inputs)
//  syndrom[ 5]:  x   x x     xx   x  (6 inputs)
//  syndrom[ 6]:   xx     x     x  xx (6 inputs)
//  syndrom[ 7]:   xx     xxxx        (6 inputs)
//  syndrom[ 8]:   x x   x  x   x x   (6 inputs)
//  syndrom[ 9]:    xx   x  x   xx    (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 6 7 9)
//  input bit  4 used  3 times (syndrom bits 3 8 9)
//  input bit  5 used  3 times (syndrom bits 0 4 5)
//  input bit  6 used  3 times (syndrom bits 1 2 4)
//  input bit  7 used  3 times (syndrom bits 1 2 5)
//  input bit  8 used  3 times (syndrom bits 0 8 9)
//  input bit  9 used  3 times (syndrom bits 3 6 7)
//  input bit 10 used  3 times (syndrom bits 0 3 7)
//  input bit 11 used  3 times (syndrom bits 7 8 9)
//  input bit 12 used  3 times (syndrom bits 1 2 7)
//  input bit 13 used  3 times (syndrom bits 1 4 5)
//  input bit 14 used  3 times (syndrom bits 2 4 5)
//  input bit 15 used  3 times (syndrom bits 6 8 9)
//  input bit 16 used  3 times (syndrom bits 0 3 9)
//  input bit 17 used  3 times (syndrom bits 0 3 8)
//  input bit 18 used  3 times (syndrom bits 4 5 6)
//  input bit 19 used  3 times (syndrom bits 1 2 6)
function [10-1:0] extended_hamming_code_30_20_f;
    input [20-1:0] in;
    reg [10-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 5]^in[ 8]^in[10]^in[16]^in[17];//6 inputs
        syndrom[ 1] = in[ 0]^in[ 6]^in[ 7]^in[12]^in[13]^in[19];//6 inputs
        syndrom[ 2] = in[ 0]^in[ 6]^in[ 7]^in[12]^in[14]^in[19];//6 inputs
        syndrom[ 3] = in[ 1]^in[ 4]^in[ 9]^in[10]^in[16]^in[17];//6 inputs
        syndrom[ 4] = in[ 1]^in[ 5]^in[ 6]^in[13]^in[14]^in[18];//6 inputs
        syndrom[ 5] = in[ 1]^in[ 5]^in[ 7]^in[13]^in[14]^in[18];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 3]^in[ 9]^in[15]^in[18]^in[19];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 3]^in[ 9]^in[10]^in[11]^in[12];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 4]^in[ 8]^in[11]^in[15]^in[17];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 4]^in[ 8]^in[11]^in[15]^in[16];//6 inputs
        extended_hamming_code_30_20_f = syndrom;
    end
endfunction
function [2+20-1:0] extended_hamming_code_30_20_f_correction_pattern_f;
    input [10-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [20-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {20{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			10'b0000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {20{1'b0}};
			end	
			10'b0000000111: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 0]=1'b1;
			end
			10'b0000111000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 1]=1'b1;
			end
			10'b0111000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 2]=1'b1;
			end
			10'b1011000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 3]=1'b1;
			end
			10'b1100001000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 4]=1'b1;
			end
			10'b0000110001: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 5]=1'b1;
			end
			10'b0000010110: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 6]=1'b1;
			end
			10'b0000100110: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 7]=1'b1;
			end
			10'b1100000001: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 8]=1'b1;
			end
			10'b0011001000: begin
				correction_pattern = {20{1'b0}};correction_pattern[ 9]=1'b1;
			end
			10'b0010001001: begin
				correction_pattern = {20{1'b0}};correction_pattern[10]=1'b1;
			end
			10'b1110000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[11]=1'b1;
			end
			10'b0010000110: begin
				correction_pattern = {20{1'b0}};correction_pattern[12]=1'b1;
			end
			10'b0000110010: begin
				correction_pattern = {20{1'b0}};correction_pattern[13]=1'b1;
			end
			10'b0000110100: begin
				correction_pattern = {20{1'b0}};correction_pattern[14]=1'b1;
			end
			10'b1101000000: begin
				correction_pattern = {20{1'b0}};correction_pattern[15]=1'b1;
			end
			10'b1000001001: begin
				correction_pattern = {20{1'b0}};correction_pattern[16]=1'b1;
			end
			10'b0100001001: begin
				correction_pattern = {20{1'b0}};correction_pattern[17]=1'b1;
			end
			10'b0001110000: begin
				correction_pattern = {20{1'b0}};correction_pattern[18]=1'b1;
			end
			10'b0001000110: begin
				correction_pattern = {20{1'b0}};correction_pattern[19]=1'b1;
			end
			10'b0000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b0100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			10'b1000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {20{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_30_20_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [10-1:0] stored_data_edc = extended_hamming_code_30_20_f(i_stored_data);
wire [10-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [20-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_30_20_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_24_balanced (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [12-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [12-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_36_24_f
//Compute 12 bits Error Detection Code from a 24 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 68719476736 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[ 0]: x x x     x x            (5 inputs)
//  syndrom[ 1]: x          x x        x  (4 inputs)
//  syndrom[ 2]:  x        x  x         x (4 inputs)
//  syndrom[ 3]:  x         xx            (3 inputs)
//  syndrom[ 4]:         x     x      x x (4 inputs)
//  syndrom[ 5]:   x      x     x  x      (4 inputs)
//  syndrom[ 6]:    x    x      x   x     (4 inputs)
//  syndrom[ 7]:    x     x    x     x    (4 inputs)
//  syndrom[ 8]:       x         x    xx  (4 inputs)
//  syndrom[ 9]:     x  x         xx      (4 inputs)
//  syndrom[10]:      xx          x x     (4 inputs)
//  syndrom[11]:      x x        x   x    (4 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 0 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 0 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 8 10)
//  input bit  7 used  2 times (syndrom bits 9 11)
//  input bit  8 used  2 times (syndrom bits 4 6)
//  input bit  9 used  2 times (syndrom bits 5 7)
//  input bit 10 used  2 times (syndrom bits 0 2)
//  input bit 11 used  2 times (syndrom bits 1 3)
//  input bit 12 used  2 times (syndrom bits 0 3)
//  input bit 13 used  2 times (syndrom bits 1 2)
//  input bit 14 used  2 times (syndrom bits 4 7)
//  input bit 15 used  2 times (syndrom bits 5 6)
//  input bit 16 used  2 times (syndrom bits 8 11)
//  input bit 17 used  2 times (syndrom bits 9 10)
//  input bit 18 used  2 times (syndrom bits 5 9)
//  input bit 19 used  2 times (syndrom bits 6 10)
//  input bit 20 used  2 times (syndrom bits 7 11)
//  input bit 21 used  2 times (syndrom bits 4 8)
//  input bit 22 used  2 times (syndrom bits 1 8)
//  input bit 23 used  2 times (syndrom bits 2 4)
function [12-1:0] hamming_code_36_24_f;
    input [24-1:0] in;
    reg [12-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 2]^in[ 4]^in[10]^in[12];//5 inputs
        syndrom[ 1] = in[ 0]^in[11]^in[13]^in[22];//4 inputs
        syndrom[ 2] = in[ 1]^in[10]^in[13]^in[23];//4 inputs
        syndrom[ 3] = in[ 1]^in[11]^in[12];//3 inputs
        syndrom[ 4] = in[ 8]^in[14]^in[21]^in[23];//4 inputs
        syndrom[ 5] = in[ 2]^in[ 9]^in[15]^in[18];//4 inputs
        syndrom[ 6] = in[ 3]^in[ 8]^in[15]^in[19];//4 inputs
        syndrom[ 7] = in[ 3]^in[ 9]^in[14]^in[20];//4 inputs
        syndrom[ 8] = in[ 6]^in[16]^in[21]^in[22];//4 inputs
        syndrom[ 9] = in[ 4]^in[ 7]^in[17]^in[18];//4 inputs
        syndrom[10] = in[ 5]^in[ 6]^in[17]^in[19];//4 inputs
        syndrom[11] = in[ 5]^in[ 7]^in[16]^in[20];//4 inputs
        hamming_code_36_24_f = syndrom;
    end
endfunction
wire [12-1:0] stored_data_edc = hamming_code_36_24_f(i_stored_data);
wire [12-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_24_balanced (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [12-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [12-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_36_24_f
//Compute 12 bits Error Detection Code from a 24 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 68719476736 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[ 0]: x     x  x     xx     x  (6 inputs)
//  syndrom[ 1]: x      xx      xx      x (6 inputs)
//  syndrom[ 2]: x      x x    x  x    x  (6 inputs)
//  syndrom[ 3]:  x    x x      x x    x  (6 inputs)
//  syndrom[ 4]:  x    x  x    x x      x (6 inputs)
//  syndrom[ 5]:  x     xx     x  x     x (6 inputs)
//  syndrom[ 6]:   x x      x x    x x    (6 inputs)
//  syndrom[ 7]:   x  x    x  x    x  x   (6 inputs)
//  syndrom[ 8]:   x  x     xx      xx    (6 inputs)
//  syndrom[ 9]:    xx     x  x     xx    (6 inputs)
//  syndrom[10]:    xx      xx     x  x   (6 inputs)
//  syndrom[11]:    x x    x x      x x   (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 6 9 10)
//  input bit  5 used  3 times (syndrom bits 7 8 11)
//  input bit  6 used  3 times (syndrom bits 0 3 4)
//  input bit  7 used  3 times (syndrom bits 1 2 5)
//  input bit  8 used  3 times (syndrom bits 1 3 5)
//  input bit  9 used  3 times (syndrom bits 0 2 4)
//  input bit 10 used  3 times (syndrom bits 7 9 11)
//  input bit 11 used  3 times (syndrom bits 6 8 10)
//  input bit 12 used  3 times (syndrom bits 8 10 11)
//  input bit 13 used  3 times (syndrom bits 6 7 9)
//  input bit 14 used  3 times (syndrom bits 2 4 5)
//  input bit 15 used  3 times (syndrom bits 0 1 3)
//  input bit 16 used  3 times (syndrom bits 0 1 4)
//  input bit 17 used  3 times (syndrom bits 2 3 5)
//  input bit 18 used  3 times (syndrom bits 6 7 10)
//  input bit 19 used  3 times (syndrom bits 8 9 11)
//  input bit 20 used  3 times (syndrom bits 6 8 9)
//  input bit 21 used  3 times (syndrom bits 7 10 11)
//  input bit 22 used  3 times (syndrom bits 0 2 3)
//  input bit 23 used  3 times (syndrom bits 1 4 5)
function [12-1:0] extended_hamming_code_36_24_f;
    input [24-1:0] in;
    reg [12-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 6]^in[ 9]^in[15]^in[16]^in[22];//6 inputs
        syndrom[ 1] = in[ 0]^in[ 7]^in[ 8]^in[15]^in[16]^in[23];//6 inputs
        syndrom[ 2] = in[ 0]^in[ 7]^in[ 9]^in[14]^in[17]^in[22];//6 inputs
        syndrom[ 3] = in[ 1]^in[ 6]^in[ 8]^in[15]^in[17]^in[22];//6 inputs
        syndrom[ 4] = in[ 1]^in[ 6]^in[ 9]^in[14]^in[16]^in[23];//6 inputs
        syndrom[ 5] = in[ 1]^in[ 7]^in[ 8]^in[14]^in[17]^in[23];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 4]^in[11]^in[13]^in[18]^in[20];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 5]^in[10]^in[13]^in[18]^in[21];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 5]^in[11]^in[12]^in[19]^in[20];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 4]^in[10]^in[13]^in[19]^in[20];//6 inputs
        syndrom[10] = in[ 3]^in[ 4]^in[11]^in[12]^in[18]^in[21];//6 inputs
        syndrom[11] = in[ 3]^in[ 5]^in[10]^in[12]^in[19]^in[21];//6 inputs
        extended_hamming_code_36_24_f = syndrom;
    end
endfunction
wire [12-1:0] stored_data_edc = extended_hamming_code_36_24_f(i_stored_data);
wire [12-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_24_balanced (
	input wire [24-1:0] i_write_data, // Data to write to storage
	output reg [12-1:0] o_write_edc, // EDC bits to write to storage
	input wire [24-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [12-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [24-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_36_24_f
//Compute 12 bits Error Detection Code from a 24 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 16777216 valid code words out of 68719476736 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[23]
//  syndrom[ 0]: x     x  x     xx     x  (6 inputs)
//  syndrom[ 1]: x      xx      xx      x (6 inputs)
//  syndrom[ 2]: x      x x    x  x    x  (6 inputs)
//  syndrom[ 3]:  x    x x      x x    x  (6 inputs)
//  syndrom[ 4]:  x    x  x    x x      x (6 inputs)
//  syndrom[ 5]:  x     xx     x  x     x (6 inputs)
//  syndrom[ 6]:   x x      x x    x x    (6 inputs)
//  syndrom[ 7]:   x  x    x  x    x  x   (6 inputs)
//  syndrom[ 8]:   x  x     xx      xx    (6 inputs)
//  syndrom[ 9]:    xx     x  x     xx    (6 inputs)
//  syndrom[10]:    xx      xx     x  x   (6 inputs)
//  syndrom[11]:    x x    x x      x x   (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 6 9 10)
//  input bit  5 used  3 times (syndrom bits 7 8 11)
//  input bit  6 used  3 times (syndrom bits 0 3 4)
//  input bit  7 used  3 times (syndrom bits 1 2 5)
//  input bit  8 used  3 times (syndrom bits 1 3 5)
//  input bit  9 used  3 times (syndrom bits 0 2 4)
//  input bit 10 used  3 times (syndrom bits 7 9 11)
//  input bit 11 used  3 times (syndrom bits 6 8 10)
//  input bit 12 used  3 times (syndrom bits 8 10 11)
//  input bit 13 used  3 times (syndrom bits 6 7 9)
//  input bit 14 used  3 times (syndrom bits 2 4 5)
//  input bit 15 used  3 times (syndrom bits 0 1 3)
//  input bit 16 used  3 times (syndrom bits 0 1 4)
//  input bit 17 used  3 times (syndrom bits 2 3 5)
//  input bit 18 used  3 times (syndrom bits 6 7 10)
//  input bit 19 used  3 times (syndrom bits 8 9 11)
//  input bit 20 used  3 times (syndrom bits 6 8 9)
//  input bit 21 used  3 times (syndrom bits 7 10 11)
//  input bit 22 used  3 times (syndrom bits 0 2 3)
//  input bit 23 used  3 times (syndrom bits 1 4 5)
function [12-1:0] extended_hamming_code_36_24_f;
    input [24-1:0] in;
    reg [12-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 6]^in[ 9]^in[15]^in[16]^in[22];//6 inputs
        syndrom[ 1] = in[ 0]^in[ 7]^in[ 8]^in[15]^in[16]^in[23];//6 inputs
        syndrom[ 2] = in[ 0]^in[ 7]^in[ 9]^in[14]^in[17]^in[22];//6 inputs
        syndrom[ 3] = in[ 1]^in[ 6]^in[ 8]^in[15]^in[17]^in[22];//6 inputs
        syndrom[ 4] = in[ 1]^in[ 6]^in[ 9]^in[14]^in[16]^in[23];//6 inputs
        syndrom[ 5] = in[ 1]^in[ 7]^in[ 8]^in[14]^in[17]^in[23];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 4]^in[11]^in[13]^in[18]^in[20];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 5]^in[10]^in[13]^in[18]^in[21];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 5]^in[11]^in[12]^in[19]^in[20];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 4]^in[10]^in[13]^in[19]^in[20];//6 inputs
        syndrom[10] = in[ 3]^in[ 4]^in[11]^in[12]^in[18]^in[21];//6 inputs
        syndrom[11] = in[ 3]^in[ 5]^in[10]^in[12]^in[19]^in[21];//6 inputs
        extended_hamming_code_36_24_f = syndrom;
    end
endfunction
function [2+24-1:0] extended_hamming_code_36_24_f_correction_pattern_f;
    input [12-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [24-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {24{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			12'b000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {24{1'b0}};
			end	
			12'b000000000111: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 0]=1'b1;
			end
			12'b000000111000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 1]=1'b1;
			end
			12'b000111000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 2]=1'b1;
			end
			12'b111000000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 3]=1'b1;
			end
			12'b011001000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 4]=1'b1;
			end
			12'b100110000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 5]=1'b1;
			end
			12'b000000011001: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 6]=1'b1;
			end
			12'b000000100110: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 7]=1'b1;
			end
			12'b000000101010: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 8]=1'b1;
			end
			12'b000000010101: begin
				correction_pattern = {24{1'b0}};correction_pattern[ 9]=1'b1;
			end
			12'b101010000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[10]=1'b1;
			end
			12'b010101000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[11]=1'b1;
			end
			12'b110100000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[12]=1'b1;
			end
			12'b001011000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[13]=1'b1;
			end
			12'b000000110100: begin
				correction_pattern = {24{1'b0}};correction_pattern[14]=1'b1;
			end
			12'b000000001011: begin
				correction_pattern = {24{1'b0}};correction_pattern[15]=1'b1;
			end
			12'b000000010011: begin
				correction_pattern = {24{1'b0}};correction_pattern[16]=1'b1;
			end
			12'b000000101100: begin
				correction_pattern = {24{1'b0}};correction_pattern[17]=1'b1;
			end
			12'b010011000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[18]=1'b1;
			end
			12'b101100000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[19]=1'b1;
			end
			12'b001101000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[20]=1'b1;
			end
			12'b110010000000: begin
				correction_pattern = {24{1'b0}};correction_pattern[21]=1'b1;
			end
			12'b000000001101: begin
				correction_pattern = {24{1'b0}};correction_pattern[22]=1'b1;
			end
			12'b000000110010: begin
				correction_pattern = {24{1'b0}};correction_pattern[23]=1'b1;
			end
			12'b000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			12'b100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {24{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_36_24_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [12-1:0] stored_data_edc = extended_hamming_code_36_24_f(i_stored_data);
wire [12-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [24-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_36_24_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_32_balanced (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [16-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [16-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_48_32_f
//Compute 16 bits Error Detection Code from a 32 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 281474976710656 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[ 0]: x             x x              x (4 inputs)
//  syndrom[ 1]: x              x x          x    (4 inputs)
//  syndrom[ 2]:  x            x  x           x   (4 inputs)
//  syndrom[ 3]:  x             xx             x  (4 inputs)
//  syndrom[ 4]:   x         x     x            x (4 inputs)
//  syndrom[ 5]:   x          x     x        x    (4 inputs)
//  syndrom[ 6]:    x        x      x         x   (4 inputs)
//  syndrom[ 7]:    x         x    x           x  (4 inputs)
//  syndrom[ 8]:     x     x         x      x     (4 inputs)
//  syndrom[ 9]:     x      x         x  x        (4 inputs)
//  syndrom[10]:      x    x          x   x       (4 inputs)
//  syndrom[11]:      x     x        x     x      (4 inputs)
//  syndrom[12]:       x x             x    x     (4 inputs)
//  syndrom[13]:       x  x             xx        (4 inputs)
//  syndrom[14]:        xx              x x       (4 inputs)
//  syndrom[15]:        x x            x   x      (4 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 12 14)
//  input bit  9 used  2 times (syndrom bits 13 15)
//  input bit 10 used  2 times (syndrom bits 8 10)
//  input bit 11 used  2 times (syndrom bits 9 11)
//  input bit 12 used  2 times (syndrom bits 4 6)
//  input bit 13 used  2 times (syndrom bits 5 7)
//  input bit 14 used  2 times (syndrom bits 0 2)
//  input bit 15 used  2 times (syndrom bits 1 3)
//  input bit 16 used  2 times (syndrom bits 0 3)
//  input bit 17 used  2 times (syndrom bits 1 2)
//  input bit 18 used  2 times (syndrom bits 4 7)
//  input bit 19 used  2 times (syndrom bits 5 6)
//  input bit 20 used  2 times (syndrom bits 8 11)
//  input bit 21 used  2 times (syndrom bits 9 10)
//  input bit 22 used  2 times (syndrom bits 12 15)
//  input bit 23 used  2 times (syndrom bits 13 14)
//  input bit 24 used  2 times (syndrom bits 9 13)
//  input bit 25 used  2 times (syndrom bits 10 14)
//  input bit 26 used  2 times (syndrom bits 11 15)
//  input bit 27 used  2 times (syndrom bits 8 12)
//  input bit 28 used  2 times (syndrom bits 1 5)
//  input bit 29 used  2 times (syndrom bits 2 6)
//  input bit 30 used  2 times (syndrom bits 3 7)
//  input bit 31 used  2 times (syndrom bits 0 4)
function [16-1:0] hamming_code_48_32_f;
    input [32-1:0] in;
    reg [16-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[14]^in[16]^in[31];//4 inputs
        syndrom[ 1] = in[ 0]^in[15]^in[17]^in[28];//4 inputs
        syndrom[ 2] = in[ 1]^in[14]^in[17]^in[29];//4 inputs
        syndrom[ 3] = in[ 1]^in[15]^in[16]^in[30];//4 inputs
        syndrom[ 4] = in[ 2]^in[12]^in[18]^in[31];//4 inputs
        syndrom[ 5] = in[ 2]^in[13]^in[19]^in[28];//4 inputs
        syndrom[ 6] = in[ 3]^in[12]^in[19]^in[29];//4 inputs
        syndrom[ 7] = in[ 3]^in[13]^in[18]^in[30];//4 inputs
        syndrom[ 8] = in[ 4]^in[10]^in[20]^in[27];//4 inputs
        syndrom[ 9] = in[ 4]^in[11]^in[21]^in[24];//4 inputs
        syndrom[10] = in[ 5]^in[10]^in[21]^in[25];//4 inputs
        syndrom[11] = in[ 5]^in[11]^in[20]^in[26];//4 inputs
        syndrom[12] = in[ 6]^in[ 8]^in[22]^in[27];//4 inputs
        syndrom[13] = in[ 6]^in[ 9]^in[23]^in[24];//4 inputs
        syndrom[14] = in[ 7]^in[ 8]^in[23]^in[25];//4 inputs
        syndrom[15] = in[ 7]^in[ 9]^in[22]^in[26];//4 inputs
        hamming_code_48_32_f = syndrom;
    end
endfunction
wire [16-1:0] stored_data_edc = hamming_code_48_32_f(i_stored_data);
wire [16-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_32_balanced (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [16-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [16-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_48_32_f
//Compute 16 bits Error Detection Code from a 32 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 281474976710656 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[ 0]: x        x  x     x     x   x    (6 inputs)
//  syndrom[ 1]: x         xx        xx         x (6 inputs)
//  syndrom[ 2]: x         xx        x x        x (6 inputs)
//  syndrom[ 3]:  x      x    x    x     x   x    (6 inputs)
//  syndrom[ 4]:  x       xx          xx       x  (6 inputs)
//  syndrom[ 5]:  x       x x         xx       x  (6 inputs)
//  syndrom[ 6]:   x    x      x x         xx     (6 inputs)
//  syndrom[ 7]:   x     x   x      x   x     x   (6 inputs)
//  syndrom[ 8]:   x     x   x      x   x     x   (6 inputs)
//  syndrom[ 9]:    x  x        xx         xx     (6 inputs)
//  syndrom[10]:    x   x     x         x      xx (6 inputs)
//  syndrom[11]:    x   x     x    xxx            (6 inputs)
//  syndrom[12]:     xx         xx        x  x    (6 inputs)
//  syndrom[13]:     xx         x x      x    x   (6 inputs)
//  syndrom[14]:     x x       x  x       x x     (6 inputs)
//  syndrom[15]:      xx       x  x       xx      (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 12 13 15)
//  input bit  6 used  3 times (syndrom bits 9 14 15)
//  input bit  7 used  3 times (syndrom bits 6 10 11)
//  input bit  8 used  3 times (syndrom bits 3 7 8)
//  input bit  9 used  3 times (syndrom bits 0 4 5)
//  input bit 10 used  3 times (syndrom bits 1 2 4)
//  input bit 11 used  3 times (syndrom bits 1 2 5)
//  input bit 12 used  3 times (syndrom bits 0 7 8)
//  input bit 13 used  3 times (syndrom bits 3 10 11)
//  input bit 14 used  3 times (syndrom bits 6 14 15)
//  input bit 15 used  3 times (syndrom bits 9 12 13)
//  input bit 16 used  3 times (syndrom bits 6 9 12)
//  input bit 17 used  3 times (syndrom bits 13 14 15)
//  input bit 18 used  3 times (syndrom bits 0 3 11)
//  input bit 19 used  3 times (syndrom bits 7 8 11)
//  input bit 20 used  3 times (syndrom bits 1 2 11)
//  input bit 21 used  3 times (syndrom bits 1 4 5)
//  input bit 22 used  3 times (syndrom bits 2 4 5)
//  input bit 23 used  3 times (syndrom bits 7 8 10)
//  input bit 24 used  3 times (syndrom bits 0 3 13)
//  input bit 25 used  3 times (syndrom bits 12 14 15)
//  input bit 26 used  3 times (syndrom bits 6 9 15)
//  input bit 27 used  3 times (syndrom bits 6 9 14)
//  input bit 28 used  3 times (syndrom bits 0 3 12)
//  input bit 29 used  3 times (syndrom bits 7 8 13)
//  input bit 30 used  3 times (syndrom bits 4 5 10)
//  input bit 31 used  3 times (syndrom bits 1 2 10)
function [16-1:0] extended_hamming_code_48_32_f;
    input [32-1:0] in;
    reg [16-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 9]^in[12]^in[18]^in[24]^in[28];//6 inputs
        syndrom[ 1] = in[ 0]^in[10]^in[11]^in[20]^in[21]^in[31];//6 inputs
        syndrom[ 2] = in[ 0]^in[10]^in[11]^in[20]^in[22]^in[31];//6 inputs
        syndrom[ 3] = in[ 1]^in[ 8]^in[13]^in[18]^in[24]^in[28];//6 inputs
        syndrom[ 4] = in[ 1]^in[ 9]^in[10]^in[21]^in[22]^in[30];//6 inputs
        syndrom[ 5] = in[ 1]^in[ 9]^in[11]^in[21]^in[22]^in[30];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 7]^in[14]^in[16]^in[26]^in[27];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 8]^in[12]^in[19]^in[23]^in[29];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 8]^in[12]^in[19]^in[23]^in[29];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 6]^in[15]^in[16]^in[26]^in[27];//6 inputs
        syndrom[10] = in[ 3]^in[ 7]^in[13]^in[23]^in[30]^in[31];//6 inputs
        syndrom[11] = in[ 3]^in[ 7]^in[13]^in[18]^in[19]^in[20];//6 inputs
        syndrom[12] = in[ 4]^in[ 5]^in[15]^in[16]^in[25]^in[28];//6 inputs
        syndrom[13] = in[ 4]^in[ 5]^in[15]^in[17]^in[24]^in[29];//6 inputs
        syndrom[14] = in[ 4]^in[ 6]^in[14]^in[17]^in[25]^in[27];//6 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[14]^in[17]^in[25]^in[26];//6 inputs
        extended_hamming_code_48_32_f = syndrom;
    end
endfunction
wire [16-1:0] stored_data_edc = extended_hamming_code_48_32_f(i_stored_data);
wire [16-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_32_balanced (
	input wire [32-1:0] i_write_data, // Data to write to storage
	output reg [16-1:0] o_write_edc, // EDC bits to write to storage
	input wire [32-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [16-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [32-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_48_32_f
//Compute 16 bits Error Detection Code from a 32 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 4294967296 valid code words out of 281474976710656 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[31]
//  syndrom[ 0]: x        x  x     x     x   x    (6 inputs)
//  syndrom[ 1]: x         xx        xx         x (6 inputs)
//  syndrom[ 2]: x         xx        x x        x (6 inputs)
//  syndrom[ 3]:  x      x    x    x     x   x    (6 inputs)
//  syndrom[ 4]:  x       xx          xx       x  (6 inputs)
//  syndrom[ 5]:  x       x x         xx       x  (6 inputs)
//  syndrom[ 6]:   x    x      x x         xx     (6 inputs)
//  syndrom[ 7]:   x     x   x      x   x     x   (6 inputs)
//  syndrom[ 8]:   x     x   x      x   x     x   (6 inputs)
//  syndrom[ 9]:    x  x        xx         xx     (6 inputs)
//  syndrom[10]:    x   x     x         x      xx (6 inputs)
//  syndrom[11]:    x   x     x    xxx            (6 inputs)
//  syndrom[12]:     xx         xx        x  x    (6 inputs)
//  syndrom[13]:     xx         x x      x    x   (6 inputs)
//  syndrom[14]:     x x       x  x       x x     (6 inputs)
//  syndrom[15]:      xx       x  x       xx      (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 12 13 15)
//  input bit  6 used  3 times (syndrom bits 9 14 15)
//  input bit  7 used  3 times (syndrom bits 6 10 11)
//  input bit  8 used  3 times (syndrom bits 3 7 8)
//  input bit  9 used  3 times (syndrom bits 0 4 5)
//  input bit 10 used  3 times (syndrom bits 1 2 4)
//  input bit 11 used  3 times (syndrom bits 1 2 5)
//  input bit 12 used  3 times (syndrom bits 0 7 8)
//  input bit 13 used  3 times (syndrom bits 3 10 11)
//  input bit 14 used  3 times (syndrom bits 6 14 15)
//  input bit 15 used  3 times (syndrom bits 9 12 13)
//  input bit 16 used  3 times (syndrom bits 6 9 12)
//  input bit 17 used  3 times (syndrom bits 13 14 15)
//  input bit 18 used  3 times (syndrom bits 0 3 11)
//  input bit 19 used  3 times (syndrom bits 7 8 11)
//  input bit 20 used  3 times (syndrom bits 1 2 11)
//  input bit 21 used  3 times (syndrom bits 1 4 5)
//  input bit 22 used  3 times (syndrom bits 2 4 5)
//  input bit 23 used  3 times (syndrom bits 7 8 10)
//  input bit 24 used  3 times (syndrom bits 0 3 13)
//  input bit 25 used  3 times (syndrom bits 12 14 15)
//  input bit 26 used  3 times (syndrom bits 6 9 15)
//  input bit 27 used  3 times (syndrom bits 6 9 14)
//  input bit 28 used  3 times (syndrom bits 0 3 12)
//  input bit 29 used  3 times (syndrom bits 7 8 13)
//  input bit 30 used  3 times (syndrom bits 4 5 10)
//  input bit 31 used  3 times (syndrom bits 1 2 10)
function [16-1:0] extended_hamming_code_48_32_f;
    input [32-1:0] in;
    reg [16-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 9]^in[12]^in[18]^in[24]^in[28];//6 inputs
        syndrom[ 1] = in[ 0]^in[10]^in[11]^in[20]^in[21]^in[31];//6 inputs
        syndrom[ 2] = in[ 0]^in[10]^in[11]^in[20]^in[22]^in[31];//6 inputs
        syndrom[ 3] = in[ 1]^in[ 8]^in[13]^in[18]^in[24]^in[28];//6 inputs
        syndrom[ 4] = in[ 1]^in[ 9]^in[10]^in[21]^in[22]^in[30];//6 inputs
        syndrom[ 5] = in[ 1]^in[ 9]^in[11]^in[21]^in[22]^in[30];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 7]^in[14]^in[16]^in[26]^in[27];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 8]^in[12]^in[19]^in[23]^in[29];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 8]^in[12]^in[19]^in[23]^in[29];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 6]^in[15]^in[16]^in[26]^in[27];//6 inputs
        syndrom[10] = in[ 3]^in[ 7]^in[13]^in[23]^in[30]^in[31];//6 inputs
        syndrom[11] = in[ 3]^in[ 7]^in[13]^in[18]^in[19]^in[20];//6 inputs
        syndrom[12] = in[ 4]^in[ 5]^in[15]^in[16]^in[25]^in[28];//6 inputs
        syndrom[13] = in[ 4]^in[ 5]^in[15]^in[17]^in[24]^in[29];//6 inputs
        syndrom[14] = in[ 4]^in[ 6]^in[14]^in[17]^in[25]^in[27];//6 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[14]^in[17]^in[25]^in[26];//6 inputs
        extended_hamming_code_48_32_f = syndrom;
    end
endfunction
function [2+32-1:0] extended_hamming_code_48_32_f_correction_pattern_f;
    input [16-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [32-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {32{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			16'b0000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {32{1'b0}};
			end	
			16'b0000000000000111: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 0]=1'b1;
			end
			16'b0000000000111000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 1]=1'b1;
			end
			16'b0000000111000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 2]=1'b1;
			end
			16'b0000111000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 3]=1'b1;
			end
			16'b0111000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 4]=1'b1;
			end
			16'b1011000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 5]=1'b1;
			end
			16'b1100001000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 6]=1'b1;
			end
			16'b0000110001000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 7]=1'b1;
			end
			16'b0000000110001000: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 8]=1'b1;
			end
			16'b0000000000110001: begin
				correction_pattern = {32{1'b0}};correction_pattern[ 9]=1'b1;
			end
			16'b0000000000010110: begin
				correction_pattern = {32{1'b0}};correction_pattern[10]=1'b1;
			end
			16'b0000000000100110: begin
				correction_pattern = {32{1'b0}};correction_pattern[11]=1'b1;
			end
			16'b0000000110000001: begin
				correction_pattern = {32{1'b0}};correction_pattern[12]=1'b1;
			end
			16'b0000110000001000: begin
				correction_pattern = {32{1'b0}};correction_pattern[13]=1'b1;
			end
			16'b1100000001000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[14]=1'b1;
			end
			16'b0011001000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[15]=1'b1;
			end
			16'b0001001001000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[16]=1'b1;
			end
			16'b1110000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[17]=1'b1;
			end
			16'b0000100000001001: begin
				correction_pattern = {32{1'b0}};correction_pattern[18]=1'b1;
			end
			16'b0000100110000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[19]=1'b1;
			end
			16'b0000100000000110: begin
				correction_pattern = {32{1'b0}};correction_pattern[20]=1'b1;
			end
			16'b0000000000110010: begin
				correction_pattern = {32{1'b0}};correction_pattern[21]=1'b1;
			end
			16'b0000000000110100: begin
				correction_pattern = {32{1'b0}};correction_pattern[22]=1'b1;
			end
			16'b0000010110000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[23]=1'b1;
			end
			16'b0010000000001001: begin
				correction_pattern = {32{1'b0}};correction_pattern[24]=1'b1;
			end
			16'b1101000000000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[25]=1'b1;
			end
			16'b1000001001000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[26]=1'b1;
			end
			16'b0100001001000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[27]=1'b1;
			end
			16'b0001000000001001: begin
				correction_pattern = {32{1'b0}};correction_pattern[28]=1'b1;
			end
			16'b0010000110000000: begin
				correction_pattern = {32{1'b0}};correction_pattern[29]=1'b1;
			end
			16'b0000010000110000: begin
				correction_pattern = {32{1'b0}};correction_pattern[30]=1'b1;
			end
			16'b0000010000000110: begin
				correction_pattern = {32{1'b0}};correction_pattern[31]=1'b1;
			end
			16'b0000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b0100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			16'b1000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {32{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_48_32_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [16-1:0] stored_data_edc = extended_hamming_code_48_32_f(i_stored_data);
wire [16-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [32-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_48_32_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_36_balanced (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [18-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [18-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_54_36_f
//Compute 18 bits Error Detection Code from a 36 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 18014398509481984 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[ 0]: x                x  x          x     (4 inputs)
//  syndrom[ 1]: x                 xx             x   (4 inputs)
//  syndrom[ 2]:  x             x    x           x    (4 inputs)
//  syndrom[ 3]:  x              x x                x (4 inputs)
//  syndrom[ 4]:   x            x   x              x  (4 inputs)
//  syndrom[ 5]:   xx            xx                   (4 inputs)
//  syndrom[ 6]:              x       x            xx (4 inputs)
//  syndrom[ 7]:    x          x       x        x     (4 inputs)
//  syndrom[ 8]:     x        x        x         x    (4 inputs)
//  syndrom[ 9]:     x         x      x           x   (4 inputs)
//  syndrom[10]:      x     x           x      x      (4 inputs)
//  syndrom[11]:      x      x           x  x         (4 inputs)
//  syndrom[12]:       x    x            x   x        (4 inputs)
//  syndrom[13]:       x     x          x     x       (4 inputs)
//  syndrom[14]:        x x               x    x      (4 inputs)
//  syndrom[15]:        x  x               xx         (4 inputs)
//  syndrom[16]:         xx                x x        (4 inputs)
//  syndrom[17]:         x x              x   x       (4 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 5 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 14 16)
//  input bit 10 used  2 times (syndrom bits 15 17)
//  input bit 11 used  2 times (syndrom bits 10 12)
//  input bit 12 used  2 times (syndrom bits 11 13)
//  input bit 13 used  2 times (syndrom bits 6 8)
//  input bit 14 used  2 times (syndrom bits 7 9)
//  input bit 15 used  2 times (syndrom bits 2 4)
//  input bit 16 used  2 times (syndrom bits 3 5)
//  input bit 17 used  2 times (syndrom bits 0 5)
//  input bit 18 used  2 times (syndrom bits 1 3)
//  input bit 19 used  2 times (syndrom bits 1 4)
//  input bit 20 used  2 times (syndrom bits 0 2)
//  input bit 21 used  2 times (syndrom bits 6 9)
//  input bit 22 used  2 times (syndrom bits 7 8)
//  input bit 23 used  2 times (syndrom bits 10 13)
//  input bit 24 used  2 times (syndrom bits 11 12)
//  input bit 25 used  2 times (syndrom bits 14 17)
//  input bit 26 used  2 times (syndrom bits 15 16)
//  input bit 27 used  2 times (syndrom bits 11 15)
//  input bit 28 used  2 times (syndrom bits 12 16)
//  input bit 29 used  2 times (syndrom bits 13 17)
//  input bit 30 used  2 times (syndrom bits 10 14)
//  input bit 31 used  2 times (syndrom bits 0 7)
//  input bit 32 used  2 times (syndrom bits 2 8)
//  input bit 33 used  2 times (syndrom bits 1 9)
//  input bit 34 used  2 times (syndrom bits 4 6)
//  input bit 35 used  2 times (syndrom bits 3 6)
function [18-1:0] hamming_code_54_36_f;
    input [36-1:0] in;
    reg [18-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[17]^in[20]^in[31];//4 inputs
        syndrom[ 1] = in[ 0]^in[18]^in[19]^in[33];//4 inputs
        syndrom[ 2] = in[ 1]^in[15]^in[20]^in[32];//4 inputs
        syndrom[ 3] = in[ 1]^in[16]^in[18]^in[35];//4 inputs
        syndrom[ 4] = in[ 2]^in[15]^in[19]^in[34];//4 inputs
        syndrom[ 5] = in[ 2]^in[ 3]^in[16]^in[17];//4 inputs
        syndrom[ 6] = in[13]^in[21]^in[34]^in[35];//4 inputs
        syndrom[ 7] = in[ 3]^in[14]^in[22]^in[31];//4 inputs
        syndrom[ 8] = in[ 4]^in[13]^in[22]^in[32];//4 inputs
        syndrom[ 9] = in[ 4]^in[14]^in[21]^in[33];//4 inputs
        syndrom[10] = in[ 5]^in[11]^in[23]^in[30];//4 inputs
        syndrom[11] = in[ 5]^in[12]^in[24]^in[27];//4 inputs
        syndrom[12] = in[ 6]^in[11]^in[24]^in[28];//4 inputs
        syndrom[13] = in[ 6]^in[12]^in[23]^in[29];//4 inputs
        syndrom[14] = in[ 7]^in[ 9]^in[25]^in[30];//4 inputs
        syndrom[15] = in[ 7]^in[10]^in[26]^in[27];//4 inputs
        syndrom[16] = in[ 8]^in[ 9]^in[26]^in[28];//4 inputs
        syndrom[17] = in[ 8]^in[10]^in[25]^in[29];//4 inputs
        hamming_code_54_36_f = syndrom;
    end
endfunction
wire [18-1:0] stored_data_edc = hamming_code_54_36_f(i_stored_data);
wire [18-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_36_balanced (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [18-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [18-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_54_36_f
//Compute 18 bits Error Detection Code from a 36 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 18014398509481984 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[ 0]: x         x  x         xx         x  (6 inputs)
//  syndrom[ 1]: x          xx          xx          x (6 inputs)
//  syndrom[ 2]: x          x x        x  x        x  (6 inputs)
//  syndrom[ 3]:  x        x x          x x        x  (6 inputs)
//  syndrom[ 4]:  x        x  x        x x          x (6 inputs)
//  syndrom[ 5]:  x         xx         x  x         x (6 inputs)
//  syndrom[ 6]:   x     x      x     x    x     x    (6 inputs)
//  syndrom[ 7]:   x      x    x      x    x      x   (6 inputs)
//  syndrom[ 8]:   x      x     x    x      x    x    (6 inputs)
//  syndrom[ 9]:    x    x     x      x     x    x    (6 inputs)
//  syndrom[10]:    x    x      x    x     x      x   (6 inputs)
//  syndrom[11]:    x     x    x     x      x     x   (6 inputs)
//  syndrom[12]:     x x          x x        x x      (6 inputs)
//  syndrom[13]:     x  x        x  x        x  x     (6 inputs)
//  syndrom[14]:     x  x         xx          xx      (6 inputs)
//  syndrom[15]:      xx         x  x         xx      (6 inputs)
//  syndrom[16]:      xx          xx         x  x     (6 inputs)
//  syndrom[17]:      x x        x x          x x     (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 12 15 16)
//  input bit  7 used  3 times (syndrom bits 13 14 17)
//  input bit  8 used  3 times (syndrom bits 6 9 10)
//  input bit  9 used  3 times (syndrom bits 7 8 11)
//  input bit 10 used  3 times (syndrom bits 0 3 4)
//  input bit 11 used  3 times (syndrom bits 1 2 5)
//  input bit 12 used  3 times (syndrom bits 1 3 5)
//  input bit 13 used  3 times (syndrom bits 0 2 4)
//  input bit 14 used  3 times (syndrom bits 7 9 11)
//  input bit 15 used  3 times (syndrom bits 6 8 10)
//  input bit 16 used  3 times (syndrom bits 13 15 17)
//  input bit 17 used  3 times (syndrom bits 12 14 16)
//  input bit 18 used  3 times (syndrom bits 14 16 17)
//  input bit 19 used  3 times (syndrom bits 12 13 15)
//  input bit 20 used  3 times (syndrom bits 8 10 11)
//  input bit 21 used  3 times (syndrom bits 6 7 9)
//  input bit 22 used  3 times (syndrom bits 2 4 5)
//  input bit 23 used  3 times (syndrom bits 0 1 3)
//  input bit 24 used  3 times (syndrom bits 0 1 4)
//  input bit 25 used  3 times (syndrom bits 2 3 5)
//  input bit 26 used  3 times (syndrom bits 6 7 10)
//  input bit 27 used  3 times (syndrom bits 8 9 11)
//  input bit 28 used  3 times (syndrom bits 12 13 16)
//  input bit 29 used  3 times (syndrom bits 14 15 17)
//  input bit 30 used  3 times (syndrom bits 12 14 15)
//  input bit 31 used  3 times (syndrom bits 13 16 17)
//  input bit 32 used  3 times (syndrom bits 6 8 9)
//  input bit 33 used  3 times (syndrom bits 7 10 11)
//  input bit 34 used  3 times (syndrom bits 0 2 3)
//  input bit 35 used  3 times (syndrom bits 1 4 5)
function [18-1:0] extended_hamming_code_54_36_f;
    input [36-1:0] in;
    reg [18-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[10]^in[13]^in[23]^in[24]^in[34];//6 inputs
        syndrom[ 1] = in[ 0]^in[11]^in[12]^in[23]^in[24]^in[35];//6 inputs
        syndrom[ 2] = in[ 0]^in[11]^in[13]^in[22]^in[25]^in[34];//6 inputs
        syndrom[ 3] = in[ 1]^in[10]^in[12]^in[23]^in[25]^in[34];//6 inputs
        syndrom[ 4] = in[ 1]^in[10]^in[13]^in[22]^in[24]^in[35];//6 inputs
        syndrom[ 5] = in[ 1]^in[11]^in[12]^in[22]^in[25]^in[35];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 8]^in[15]^in[21]^in[26]^in[32];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 9]^in[14]^in[21]^in[26]^in[33];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 9]^in[15]^in[20]^in[27]^in[32];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 8]^in[14]^in[21]^in[27]^in[32];//6 inputs
        syndrom[10] = in[ 3]^in[ 8]^in[15]^in[20]^in[26]^in[33];//6 inputs
        syndrom[11] = in[ 3]^in[ 9]^in[14]^in[20]^in[27]^in[33];//6 inputs
        syndrom[12] = in[ 4]^in[ 6]^in[17]^in[19]^in[28]^in[30];//6 inputs
        syndrom[13] = in[ 4]^in[ 7]^in[16]^in[19]^in[28]^in[31];//6 inputs
        syndrom[14] = in[ 4]^in[ 7]^in[17]^in[18]^in[29]^in[30];//6 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[16]^in[19]^in[29]^in[30];//6 inputs
        syndrom[16] = in[ 5]^in[ 6]^in[17]^in[18]^in[28]^in[31];//6 inputs
        syndrom[17] = in[ 5]^in[ 7]^in[16]^in[18]^in[29]^in[31];//6 inputs
        extended_hamming_code_54_36_f = syndrom;
    end
endfunction
wire [18-1:0] stored_data_edc = extended_hamming_code_54_36_f(i_stored_data);
wire [18-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_36_balanced (
	input wire [36-1:0] i_write_data, // Data to write to storage
	output reg [18-1:0] o_write_edc, // EDC bits to write to storage
	input wire [36-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [18-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [36-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_54_36_f
//Compute 18 bits Error Detection Code from a 36 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 68719476736 valid code words out of 18014398509481984 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[35]
//  syndrom[ 0]: x         x  x         xx         x  (6 inputs)
//  syndrom[ 1]: x          xx          xx          x (6 inputs)
//  syndrom[ 2]: x          x x        x  x        x  (6 inputs)
//  syndrom[ 3]:  x        x x          x x        x  (6 inputs)
//  syndrom[ 4]:  x        x  x        x x          x (6 inputs)
//  syndrom[ 5]:  x         xx         x  x         x (6 inputs)
//  syndrom[ 6]:   x     x      x     x    x     x    (6 inputs)
//  syndrom[ 7]:   x      x    x      x    x      x   (6 inputs)
//  syndrom[ 8]:   x      x     x    x      x    x    (6 inputs)
//  syndrom[ 9]:    x    x     x      x     x    x    (6 inputs)
//  syndrom[10]:    x    x      x    x     x      x   (6 inputs)
//  syndrom[11]:    x     x    x     x      x     x   (6 inputs)
//  syndrom[12]:     x x          x x        x x      (6 inputs)
//  syndrom[13]:     x  x        x  x        x  x     (6 inputs)
//  syndrom[14]:     x  x         xx          xx      (6 inputs)
//  syndrom[15]:      xx         x  x         xx      (6 inputs)
//  syndrom[16]:      xx          xx         x  x     (6 inputs)
//  syndrom[17]:      x x        x x          x x     (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 12 15 16)
//  input bit  7 used  3 times (syndrom bits 13 14 17)
//  input bit  8 used  3 times (syndrom bits 6 9 10)
//  input bit  9 used  3 times (syndrom bits 7 8 11)
//  input bit 10 used  3 times (syndrom bits 0 3 4)
//  input bit 11 used  3 times (syndrom bits 1 2 5)
//  input bit 12 used  3 times (syndrom bits 1 3 5)
//  input bit 13 used  3 times (syndrom bits 0 2 4)
//  input bit 14 used  3 times (syndrom bits 7 9 11)
//  input bit 15 used  3 times (syndrom bits 6 8 10)
//  input bit 16 used  3 times (syndrom bits 13 15 17)
//  input bit 17 used  3 times (syndrom bits 12 14 16)
//  input bit 18 used  3 times (syndrom bits 14 16 17)
//  input bit 19 used  3 times (syndrom bits 12 13 15)
//  input bit 20 used  3 times (syndrom bits 8 10 11)
//  input bit 21 used  3 times (syndrom bits 6 7 9)
//  input bit 22 used  3 times (syndrom bits 2 4 5)
//  input bit 23 used  3 times (syndrom bits 0 1 3)
//  input bit 24 used  3 times (syndrom bits 0 1 4)
//  input bit 25 used  3 times (syndrom bits 2 3 5)
//  input bit 26 used  3 times (syndrom bits 6 7 10)
//  input bit 27 used  3 times (syndrom bits 8 9 11)
//  input bit 28 used  3 times (syndrom bits 12 13 16)
//  input bit 29 used  3 times (syndrom bits 14 15 17)
//  input bit 30 used  3 times (syndrom bits 12 14 15)
//  input bit 31 used  3 times (syndrom bits 13 16 17)
//  input bit 32 used  3 times (syndrom bits 6 8 9)
//  input bit 33 used  3 times (syndrom bits 7 10 11)
//  input bit 34 used  3 times (syndrom bits 0 2 3)
//  input bit 35 used  3 times (syndrom bits 1 4 5)
function [18-1:0] extended_hamming_code_54_36_f;
    input [36-1:0] in;
    reg [18-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[10]^in[13]^in[23]^in[24]^in[34];//6 inputs
        syndrom[ 1] = in[ 0]^in[11]^in[12]^in[23]^in[24]^in[35];//6 inputs
        syndrom[ 2] = in[ 0]^in[11]^in[13]^in[22]^in[25]^in[34];//6 inputs
        syndrom[ 3] = in[ 1]^in[10]^in[12]^in[23]^in[25]^in[34];//6 inputs
        syndrom[ 4] = in[ 1]^in[10]^in[13]^in[22]^in[24]^in[35];//6 inputs
        syndrom[ 5] = in[ 1]^in[11]^in[12]^in[22]^in[25]^in[35];//6 inputs
        syndrom[ 6] = in[ 2]^in[ 8]^in[15]^in[21]^in[26]^in[32];//6 inputs
        syndrom[ 7] = in[ 2]^in[ 9]^in[14]^in[21]^in[26]^in[33];//6 inputs
        syndrom[ 8] = in[ 2]^in[ 9]^in[15]^in[20]^in[27]^in[32];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 8]^in[14]^in[21]^in[27]^in[32];//6 inputs
        syndrom[10] = in[ 3]^in[ 8]^in[15]^in[20]^in[26]^in[33];//6 inputs
        syndrom[11] = in[ 3]^in[ 9]^in[14]^in[20]^in[27]^in[33];//6 inputs
        syndrom[12] = in[ 4]^in[ 6]^in[17]^in[19]^in[28]^in[30];//6 inputs
        syndrom[13] = in[ 4]^in[ 7]^in[16]^in[19]^in[28]^in[31];//6 inputs
        syndrom[14] = in[ 4]^in[ 7]^in[17]^in[18]^in[29]^in[30];//6 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[16]^in[19]^in[29]^in[30];//6 inputs
        syndrom[16] = in[ 5]^in[ 6]^in[17]^in[18]^in[28]^in[31];//6 inputs
        syndrom[17] = in[ 5]^in[ 7]^in[16]^in[18]^in[29]^in[31];//6 inputs
        extended_hamming_code_54_36_f = syndrom;
    end
endfunction
function [2+36-1:0] extended_hamming_code_54_36_f_correction_pattern_f;
    input [18-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [36-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {36{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			18'b000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {36{1'b0}};
			end	
			18'b000000000000000111: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 0]=1'b1;
			end
			18'b000000000000111000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 1]=1'b1;
			end
			18'b000000000111000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 2]=1'b1;
			end
			18'b000000111000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 3]=1'b1;
			end
			18'b000111000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 4]=1'b1;
			end
			18'b111000000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 5]=1'b1;
			end
			18'b011001000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 6]=1'b1;
			end
			18'b100110000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 7]=1'b1;
			end
			18'b000000011001000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 8]=1'b1;
			end
			18'b000000100110000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[ 9]=1'b1;
			end
			18'b000000000000011001: begin
				correction_pattern = {36{1'b0}};correction_pattern[10]=1'b1;
			end
			18'b000000000000100110: begin
				correction_pattern = {36{1'b0}};correction_pattern[11]=1'b1;
			end
			18'b000000000000101010: begin
				correction_pattern = {36{1'b0}};correction_pattern[12]=1'b1;
			end
			18'b000000000000010101: begin
				correction_pattern = {36{1'b0}};correction_pattern[13]=1'b1;
			end
			18'b000000101010000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[14]=1'b1;
			end
			18'b000000010101000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[15]=1'b1;
			end
			18'b101010000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[16]=1'b1;
			end
			18'b010101000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[17]=1'b1;
			end
			18'b110100000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[18]=1'b1;
			end
			18'b001011000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[19]=1'b1;
			end
			18'b000000110100000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[20]=1'b1;
			end
			18'b000000001011000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[21]=1'b1;
			end
			18'b000000000000110100: begin
				correction_pattern = {36{1'b0}};correction_pattern[22]=1'b1;
			end
			18'b000000000000001011: begin
				correction_pattern = {36{1'b0}};correction_pattern[23]=1'b1;
			end
			18'b000000000000010011: begin
				correction_pattern = {36{1'b0}};correction_pattern[24]=1'b1;
			end
			18'b000000000000101100: begin
				correction_pattern = {36{1'b0}};correction_pattern[25]=1'b1;
			end
			18'b000000010011000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[26]=1'b1;
			end
			18'b000000101100000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[27]=1'b1;
			end
			18'b010011000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[28]=1'b1;
			end
			18'b101100000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[29]=1'b1;
			end
			18'b001101000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[30]=1'b1;
			end
			18'b110010000000000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[31]=1'b1;
			end
			18'b000000001101000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[32]=1'b1;
			end
			18'b000000110010000000: begin
				correction_pattern = {36{1'b0}};correction_pattern[33]=1'b1;
			end
			18'b000000000000001101: begin
				correction_pattern = {36{1'b0}};correction_pattern[34]=1'b1;
			end
			18'b000000000000110010: begin
				correction_pattern = {36{1'b0}};correction_pattern[35]=1'b1;
			end
			18'b000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			18'b100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {36{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_54_36_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [18-1:0] stored_data_edc = extended_hamming_code_54_36_f(i_stored_data);
wire [18-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [36-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_54_36_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_40_balanced (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [20-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [20-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_60_40_f
//Compute 20 bits Error Detection Code from a 40 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 1152921504606846976 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[ 0]: x x x             x x                    (5 inputs)
//  syndrom[ 1]: x                  x x                x  (4 inputs)
//  syndrom[ 2]:  x                x  x                 x (4 inputs)
//  syndrom[ 3]:  x                 xx                    (3 inputs)
//  syndrom[ 4]:                 x     x              x x (4 inputs)
//  syndrom[ 5]:   x              x     x          x      (4 inputs)
//  syndrom[ 6]:    x            x      x           x     (4 inputs)
//  syndrom[ 7]:    x             x    x             x    (4 inputs)
//  syndrom[ 8]:               x         x            xx  (4 inputs)
//  syndrom[ 9]:     x          x         x        x      (4 inputs)
//  syndrom[10]:      x        x          x         x     (4 inputs)
//  syndrom[11]:      x         x        x           x    (4 inputs)
//  syndrom[12]:       x     x             x      x       (4 inputs)
//  syndrom[13]:       x      x             x  x          (4 inputs)
//  syndrom[14]:        x    x              x   x         (4 inputs)
//  syndrom[15]:        x     x            x     x        (4 inputs)
//  syndrom[16]:         x x                 x    x       (4 inputs)
//  syndrom[17]:         x  x                 xx          (4 inputs)
//  syndrom[18]:          xx                  x x         (4 inputs)
//  syndrom[19]:          x x                x   x        (4 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 0 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 0 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 16 18)
//  input bit 11 used  2 times (syndrom bits 17 19)
//  input bit 12 used  2 times (syndrom bits 12 14)
//  input bit 13 used  2 times (syndrom bits 13 15)
//  input bit 14 used  2 times (syndrom bits 8 10)
//  input bit 15 used  2 times (syndrom bits 9 11)
//  input bit 16 used  2 times (syndrom bits 4 6)
//  input bit 17 used  2 times (syndrom bits 5 7)
//  input bit 18 used  2 times (syndrom bits 0 2)
//  input bit 19 used  2 times (syndrom bits 1 3)
//  input bit 20 used  2 times (syndrom bits 0 3)
//  input bit 21 used  2 times (syndrom bits 1 2)
//  input bit 22 used  2 times (syndrom bits 4 7)
//  input bit 23 used  2 times (syndrom bits 5 6)
//  input bit 24 used  2 times (syndrom bits 8 11)
//  input bit 25 used  2 times (syndrom bits 9 10)
//  input bit 26 used  2 times (syndrom bits 12 15)
//  input bit 27 used  2 times (syndrom bits 13 14)
//  input bit 28 used  2 times (syndrom bits 16 19)
//  input bit 29 used  2 times (syndrom bits 17 18)
//  input bit 30 used  2 times (syndrom bits 13 17)
//  input bit 31 used  2 times (syndrom bits 14 18)
//  input bit 32 used  2 times (syndrom bits 15 19)
//  input bit 33 used  2 times (syndrom bits 12 16)
//  input bit 34 used  2 times (syndrom bits 5 9)
//  input bit 35 used  2 times (syndrom bits 6 10)
//  input bit 36 used  2 times (syndrom bits 7 11)
//  input bit 37 used  2 times (syndrom bits 4 8)
//  input bit 38 used  2 times (syndrom bits 1 8)
//  input bit 39 used  2 times (syndrom bits 2 4)
function [20-1:0] hamming_code_60_40_f;
    input [40-1:0] in;
    reg [20-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[ 2]^in[ 4]^in[18]^in[20];//5 inputs
        syndrom[ 1] = in[ 0]^in[19]^in[21]^in[38];//4 inputs
        syndrom[ 2] = in[ 1]^in[18]^in[21]^in[39];//4 inputs
        syndrom[ 3] = in[ 1]^in[19]^in[20];//3 inputs
        syndrom[ 4] = in[16]^in[22]^in[37]^in[39];//4 inputs
        syndrom[ 5] = in[ 2]^in[17]^in[23]^in[34];//4 inputs
        syndrom[ 6] = in[ 3]^in[16]^in[23]^in[35];//4 inputs
        syndrom[ 7] = in[ 3]^in[17]^in[22]^in[36];//4 inputs
        syndrom[ 8] = in[14]^in[24]^in[37]^in[38];//4 inputs
        syndrom[ 9] = in[ 4]^in[15]^in[25]^in[34];//4 inputs
        syndrom[10] = in[ 5]^in[14]^in[25]^in[35];//4 inputs
        syndrom[11] = in[ 5]^in[15]^in[24]^in[36];//4 inputs
        syndrom[12] = in[ 6]^in[12]^in[26]^in[33];//4 inputs
        syndrom[13] = in[ 6]^in[13]^in[27]^in[30];//4 inputs
        syndrom[14] = in[ 7]^in[12]^in[27]^in[31];//4 inputs
        syndrom[15] = in[ 7]^in[13]^in[26]^in[32];//4 inputs
        syndrom[16] = in[ 8]^in[10]^in[28]^in[33];//4 inputs
        syndrom[17] = in[ 8]^in[11]^in[29]^in[30];//4 inputs
        syndrom[18] = in[ 9]^in[10]^in[29]^in[31];//4 inputs
        syndrom[19] = in[ 9]^in[11]^in[28]^in[32];//4 inputs
        hamming_code_60_40_f = syndrom;
    end
endfunction
wire [20-1:0] stored_data_edc = hamming_code_60_40_f(i_stored_data);
wire [20-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_40_balanced (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [20-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [20-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_60_40_f
//Compute 20 bits Error Detection Code from a 40 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 1152921504606846976 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[ 0]: x           xx            xx          x  (6 inputs)
//  syndrom[ 1]: x           x x          x  x        x   (6 inputs)
//  syndrom[ 2]: x            xx         x    x      x    (6 inputs)
//  syndrom[ 3]:  x         x   x        x   x         x  (6 inputs)
//  syndrom[ 4]:  x         x   x        x   x         x  (6 inputs)
//  syndrom[ 5]:  x          xx            xx           x (6 inputs)
//  syndrom[ 6]:   x       x     x     x       x     x    (6 inputs)
//  syndrom[ 7]:   x       x     x      x     x       x   (6 inputs)
//  syndrom[ 8]:   x        x  x          x x           x (6 inputs)
//  syndrom[ 9]:    x     x       x    x       x     x    (6 inputs)
//  syndrom[10]:    x     x       x    x        x  x      (6 inputs)
//  syndrom[11]:    x      x    x         xx            x (6 inputs)
//  syndrom[12]:     x   x         x x           xx       (6 inputs)
//  syndrom[13]:     x   x         x  x         x   x     (6 inputs)
//  syndrom[14]:     x    x      x      x      x    x     (6 inputs)
//  syndrom[15]:      xx            x x         x   x     (6 inputs)
//  syndrom[16]:      x x           xx            xx      (6 inputs)
//  syndrom[17]:      x  x        x     x     x       x   (6 inputs)
//  syndrom[18]:       xx          x  x          xx       (6 inputs)
//  syndrom[19]:       xx           xx           x x      (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 15 18 19)
//  input bit  7 used  3 times (syndrom bits 16 18 19)
//  input bit  8 used  3 times (syndrom bits 12 13 17)
//  input bit  9 used  3 times (syndrom bits 9 10 14)
//  input bit 10 used  3 times (syndrom bits 6 7 11)
//  input bit 11 used  3 times (syndrom bits 3 4 8)
//  input bit 12 used  3 times (syndrom bits 0 1 5)
//  input bit 13 used  3 times (syndrom bits 0 2 5)
//  input bit 14 used  3 times (syndrom bits 1 2 8)
//  input bit 15 used  3 times (syndrom bits 3 4 11)
//  input bit 16 used  3 times (syndrom bits 6 7 14)
//  input bit 17 used  3 times (syndrom bits 9 10 17)
//  input bit 18 used  3 times (syndrom bits 12 13 18)
//  input bit 19 used  3 times (syndrom bits 15 16 19)
//  input bit 20 used  3 times (syndrom bits 12 16 19)
//  input bit 21 used  3 times (syndrom bits 13 15 18)
//  input bit 22 used  3 times (syndrom bits 6 9 10)
//  input bit 23 used  3 times (syndrom bits 7 14 17)
//  input bit 24 used  3 times (syndrom bits 2 3 4)
//  input bit 25 used  3 times (syndrom bits 1 8 11)
//  input bit 26 used  3 times (syndrom bits 0 5 11)
//  input bit 27 used  3 times (syndrom bits 0 5 8)
//  input bit 28 used  3 times (syndrom bits 1 3 4)
//  input bit 29 used  3 times (syndrom bits 2 7 17)
//  input bit 30 used  3 times (syndrom bits 6 9 14)
//  input bit 31 used  3 times (syndrom bits 10 13 15)
//  input bit 32 used  3 times (syndrom bits 12 18 19)
//  input bit 33 used  3 times (syndrom bits 12 16 18)
//  input bit 34 used  3 times (syndrom bits 10 16 19)
//  input bit 35 used  3 times (syndrom bits 13 14 15)
//  input bit 36 used  3 times (syndrom bits 2 6 9)
//  input bit 37 used  3 times (syndrom bits 1 7 17)
//  input bit 38 used  3 times (syndrom bits 0 3 4)
//  input bit 39 used  3 times (syndrom bits 5 8 11)
function [20-1:0] extended_hamming_code_60_40_f;
    input [40-1:0] in;
    reg [20-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[12]^in[13]^in[26]^in[27]^in[38];//6 inputs
        syndrom[ 1] = in[ 0]^in[12]^in[14]^in[25]^in[28]^in[37];//6 inputs
        syndrom[ 2] = in[ 0]^in[13]^in[14]^in[24]^in[29]^in[36];//6 inputs
        syndrom[ 3] = in[ 1]^in[11]^in[15]^in[24]^in[28]^in[38];//6 inputs
        syndrom[ 4] = in[ 1]^in[11]^in[15]^in[24]^in[28]^in[38];//6 inputs
        syndrom[ 5] = in[ 1]^in[12]^in[13]^in[26]^in[27]^in[39];//6 inputs
        syndrom[ 6] = in[ 2]^in[10]^in[16]^in[22]^in[30]^in[36];//6 inputs
        syndrom[ 7] = in[ 2]^in[10]^in[16]^in[23]^in[29]^in[37];//6 inputs
        syndrom[ 8] = in[ 2]^in[11]^in[14]^in[25]^in[27]^in[39];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 9]^in[17]^in[22]^in[30]^in[36];//6 inputs
        syndrom[10] = in[ 3]^in[ 9]^in[17]^in[22]^in[31]^in[34];//6 inputs
        syndrom[11] = in[ 3]^in[10]^in[15]^in[25]^in[26]^in[39];//6 inputs
        syndrom[12] = in[ 4]^in[ 8]^in[18]^in[20]^in[32]^in[33];//6 inputs
        syndrom[13] = in[ 4]^in[ 8]^in[18]^in[21]^in[31]^in[35];//6 inputs
        syndrom[14] = in[ 4]^in[ 9]^in[16]^in[23]^in[30]^in[35];//6 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[19]^in[21]^in[31]^in[35];//6 inputs
        syndrom[16] = in[ 5]^in[ 7]^in[19]^in[20]^in[33]^in[34];//6 inputs
        syndrom[17] = in[ 5]^in[ 8]^in[17]^in[23]^in[29]^in[37];//6 inputs
        syndrom[18] = in[ 6]^in[ 7]^in[18]^in[21]^in[32]^in[33];//6 inputs
        syndrom[19] = in[ 6]^in[ 7]^in[19]^in[20]^in[32]^in[34];//6 inputs
        extended_hamming_code_60_40_f = syndrom;
    end
endfunction
wire [20-1:0] stored_data_edc = extended_hamming_code_60_40_f(i_stored_data);
wire [20-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_40_balanced (
	input wire [40-1:0] i_write_data, // Data to write to storage
	output reg [20-1:0] o_write_edc, // EDC bits to write to storage
	input wire [40-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [20-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [40-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_60_40_f
//Compute 20 bits Error Detection Code from a 40 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 1099511627776 valid code words out of 1152921504606846976 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[39]
//  syndrom[ 0]: x           xx            xx          x  (6 inputs)
//  syndrom[ 1]: x           x x          x  x        x   (6 inputs)
//  syndrom[ 2]: x            xx         x    x      x    (6 inputs)
//  syndrom[ 3]:  x         x   x        x   x         x  (6 inputs)
//  syndrom[ 4]:  x         x   x        x   x         x  (6 inputs)
//  syndrom[ 5]:  x          xx            xx           x (6 inputs)
//  syndrom[ 6]:   x       x     x     x       x     x    (6 inputs)
//  syndrom[ 7]:   x       x     x      x     x       x   (6 inputs)
//  syndrom[ 8]:   x        x  x          x x           x (6 inputs)
//  syndrom[ 9]:    x     x       x    x       x     x    (6 inputs)
//  syndrom[10]:    x     x       x    x        x  x      (6 inputs)
//  syndrom[11]:    x      x    x         xx            x (6 inputs)
//  syndrom[12]:     x   x         x x           xx       (6 inputs)
//  syndrom[13]:     x   x         x  x         x   x     (6 inputs)
//  syndrom[14]:     x    x      x      x      x    x     (6 inputs)
//  syndrom[15]:      xx            x x         x   x     (6 inputs)
//  syndrom[16]:      x x           xx            xx      (6 inputs)
//  syndrom[17]:      x  x        x     x     x       x   (6 inputs)
//  syndrom[18]:       xx          x  x          xx       (6 inputs)
//  syndrom[19]:       xx           xx           x x      (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 15 18 19)
//  input bit  7 used  3 times (syndrom bits 16 18 19)
//  input bit  8 used  3 times (syndrom bits 12 13 17)
//  input bit  9 used  3 times (syndrom bits 9 10 14)
//  input bit 10 used  3 times (syndrom bits 6 7 11)
//  input bit 11 used  3 times (syndrom bits 3 4 8)
//  input bit 12 used  3 times (syndrom bits 0 1 5)
//  input bit 13 used  3 times (syndrom bits 0 2 5)
//  input bit 14 used  3 times (syndrom bits 1 2 8)
//  input bit 15 used  3 times (syndrom bits 3 4 11)
//  input bit 16 used  3 times (syndrom bits 6 7 14)
//  input bit 17 used  3 times (syndrom bits 9 10 17)
//  input bit 18 used  3 times (syndrom bits 12 13 18)
//  input bit 19 used  3 times (syndrom bits 15 16 19)
//  input bit 20 used  3 times (syndrom bits 12 16 19)
//  input bit 21 used  3 times (syndrom bits 13 15 18)
//  input bit 22 used  3 times (syndrom bits 6 9 10)
//  input bit 23 used  3 times (syndrom bits 7 14 17)
//  input bit 24 used  3 times (syndrom bits 2 3 4)
//  input bit 25 used  3 times (syndrom bits 1 8 11)
//  input bit 26 used  3 times (syndrom bits 0 5 11)
//  input bit 27 used  3 times (syndrom bits 0 5 8)
//  input bit 28 used  3 times (syndrom bits 1 3 4)
//  input bit 29 used  3 times (syndrom bits 2 7 17)
//  input bit 30 used  3 times (syndrom bits 6 9 14)
//  input bit 31 used  3 times (syndrom bits 10 13 15)
//  input bit 32 used  3 times (syndrom bits 12 18 19)
//  input bit 33 used  3 times (syndrom bits 12 16 18)
//  input bit 34 used  3 times (syndrom bits 10 16 19)
//  input bit 35 used  3 times (syndrom bits 13 14 15)
//  input bit 36 used  3 times (syndrom bits 2 6 9)
//  input bit 37 used  3 times (syndrom bits 1 7 17)
//  input bit 38 used  3 times (syndrom bits 0 3 4)
//  input bit 39 used  3 times (syndrom bits 5 8 11)
function [20-1:0] extended_hamming_code_60_40_f;
    input [40-1:0] in;
    reg [20-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[12]^in[13]^in[26]^in[27]^in[38];//6 inputs
        syndrom[ 1] = in[ 0]^in[12]^in[14]^in[25]^in[28]^in[37];//6 inputs
        syndrom[ 2] = in[ 0]^in[13]^in[14]^in[24]^in[29]^in[36];//6 inputs
        syndrom[ 3] = in[ 1]^in[11]^in[15]^in[24]^in[28]^in[38];//6 inputs
        syndrom[ 4] = in[ 1]^in[11]^in[15]^in[24]^in[28]^in[38];//6 inputs
        syndrom[ 5] = in[ 1]^in[12]^in[13]^in[26]^in[27]^in[39];//6 inputs
        syndrom[ 6] = in[ 2]^in[10]^in[16]^in[22]^in[30]^in[36];//6 inputs
        syndrom[ 7] = in[ 2]^in[10]^in[16]^in[23]^in[29]^in[37];//6 inputs
        syndrom[ 8] = in[ 2]^in[11]^in[14]^in[25]^in[27]^in[39];//6 inputs
        syndrom[ 9] = in[ 3]^in[ 9]^in[17]^in[22]^in[30]^in[36];//6 inputs
        syndrom[10] = in[ 3]^in[ 9]^in[17]^in[22]^in[31]^in[34];//6 inputs
        syndrom[11] = in[ 3]^in[10]^in[15]^in[25]^in[26]^in[39];//6 inputs
        syndrom[12] = in[ 4]^in[ 8]^in[18]^in[20]^in[32]^in[33];//6 inputs
        syndrom[13] = in[ 4]^in[ 8]^in[18]^in[21]^in[31]^in[35];//6 inputs
        syndrom[14] = in[ 4]^in[ 9]^in[16]^in[23]^in[30]^in[35];//6 inputs
        syndrom[15] = in[ 5]^in[ 6]^in[19]^in[21]^in[31]^in[35];//6 inputs
        syndrom[16] = in[ 5]^in[ 7]^in[19]^in[20]^in[33]^in[34];//6 inputs
        syndrom[17] = in[ 5]^in[ 8]^in[17]^in[23]^in[29]^in[37];//6 inputs
        syndrom[18] = in[ 6]^in[ 7]^in[18]^in[21]^in[32]^in[33];//6 inputs
        syndrom[19] = in[ 6]^in[ 7]^in[19]^in[20]^in[32]^in[34];//6 inputs
        extended_hamming_code_60_40_f = syndrom;
    end
endfunction
function [2+40-1:0] extended_hamming_code_60_40_f_correction_pattern_f;
    input [20-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [40-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {40{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			20'b00000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {40{1'b0}};
			end	
			20'b00000000000000000111: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 0]=1'b1;
			end
			20'b00000000000000111000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 1]=1'b1;
			end
			20'b00000000000111000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 2]=1'b1;
			end
			20'b00000000111000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 3]=1'b1;
			end
			20'b00000111000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 4]=1'b1;
			end
			20'b00111000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 5]=1'b1;
			end
			20'b11001000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 6]=1'b1;
			end
			20'b11010000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 7]=1'b1;
			end
			20'b00100011000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 8]=1'b1;
			end
			20'b00000100011000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[ 9]=1'b1;
			end
			20'b00000000100011000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[10]=1'b1;
			end
			20'b00000000000100011000: begin
				correction_pattern = {40{1'b0}};correction_pattern[11]=1'b1;
			end
			20'b00000000000000100011: begin
				correction_pattern = {40{1'b0}};correction_pattern[12]=1'b1;
			end
			20'b00000000000000100101: begin
				correction_pattern = {40{1'b0}};correction_pattern[13]=1'b1;
			end
			20'b00000000000100000110: begin
				correction_pattern = {40{1'b0}};correction_pattern[14]=1'b1;
			end
			20'b00000000100000011000: begin
				correction_pattern = {40{1'b0}};correction_pattern[15]=1'b1;
			end
			20'b00000100000011000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[16]=1'b1;
			end
			20'b00100000011000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[17]=1'b1;
			end
			20'b01000011000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[18]=1'b1;
			end
			20'b10011000000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[19]=1'b1;
			end
			20'b10010001000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[20]=1'b1;
			end
			20'b01001010000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[21]=1'b1;
			end
			20'b00000000011001000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[22]=1'b1;
			end
			20'b00100100000010000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[23]=1'b1;
			end
			20'b00000000000000011100: begin
				correction_pattern = {40{1'b0}};correction_pattern[24]=1'b1;
			end
			20'b00000000100100000010: begin
				correction_pattern = {40{1'b0}};correction_pattern[25]=1'b1;
			end
			20'b00000000100000100001: begin
				correction_pattern = {40{1'b0}};correction_pattern[26]=1'b1;
			end
			20'b00000000000100100001: begin
				correction_pattern = {40{1'b0}};correction_pattern[27]=1'b1;
			end
			20'b00000000000000011010: begin
				correction_pattern = {40{1'b0}};correction_pattern[28]=1'b1;
			end
			20'b00100000000010000100: begin
				correction_pattern = {40{1'b0}};correction_pattern[29]=1'b1;
			end
			20'b00000100001001000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[30]=1'b1;
			end
			20'b00001010010000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[31]=1'b1;
			end
			20'b11000001000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[32]=1'b1;
			end
			20'b01010001000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[33]=1'b1;
			end
			20'b10010000010000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[34]=1'b1;
			end
			20'b00001110000000000000: begin
				correction_pattern = {40{1'b0}};correction_pattern[35]=1'b1;
			end
			20'b00000000001001000100: begin
				correction_pattern = {40{1'b0}};correction_pattern[36]=1'b1;
			end
			20'b00100000000010000010: begin
				correction_pattern = {40{1'b0}};correction_pattern[37]=1'b1;
			end
			20'b00000000000000011001: begin
				correction_pattern = {40{1'b0}};correction_pattern[38]=1'b1;
			end
			20'b00000000100100100000: begin
				correction_pattern = {40{1'b0}};correction_pattern[39]=1'b1;
			end
			20'b00000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b00100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b01000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			20'b10000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {40{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_60_40_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [20-1:0] stored_data_edc = extended_hamming_code_60_40_f(i_stored_data);
wire [20-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [40-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_60_40_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_48_balanced (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [24-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [24-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_72_48_f
//Compute 24 bits Error Detection Code from a 48 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[ 0]: x                     x x                      x (4 inputs)
//  syndrom[ 1]: x                      x x                  x    (4 inputs)
//  syndrom[ 2]:  x                    x  x                   x   (4 inputs)
//  syndrom[ 3]:  x                     xx                     x  (4 inputs)
//  syndrom[ 4]:   x                 x     x                    x (4 inputs)
//  syndrom[ 5]:   x                  x     x                x    (4 inputs)
//  syndrom[ 6]:    x                x      x                 x   (4 inputs)
//  syndrom[ 7]:    x                 x    x                   x  (4 inputs)
//  syndrom[ 8]:     x             x         x              x     (4 inputs)
//  syndrom[ 9]:     x              x         x          x        (4 inputs)
//  syndrom[10]:      x            x          x           x       (4 inputs)
//  syndrom[11]:      x             x        x             x      (4 inputs)
//  syndrom[12]:       x         x             x            x     (4 inputs)
//  syndrom[13]:       x          x             x        x        (4 inputs)
//  syndrom[14]:        x        x              x         x       (4 inputs)
//  syndrom[15]:        x         x            x           x      (4 inputs)
//  syndrom[16]:         x     x                 x      x         (4 inputs)
//  syndrom[17]:         x      x                 x  x            (4 inputs)
//  syndrom[18]:          x    x                  x   x           (4 inputs)
//  syndrom[19]:          x     x                x     x          (4 inputs)
//  syndrom[20]:           x x                     x    x         (4 inputs)
//  syndrom[21]:           x  x                     xx            (4 inputs)
//  syndrom[22]:            xx                      x x           (4 inputs)
//  syndrom[23]:            x x                    x   x          (4 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 20 22)
//  input bit 13 used  2 times (syndrom bits 21 23)
//  input bit 14 used  2 times (syndrom bits 16 18)
//  input bit 15 used  2 times (syndrom bits 17 19)
//  input bit 16 used  2 times (syndrom bits 12 14)
//  input bit 17 used  2 times (syndrom bits 13 15)
//  input bit 18 used  2 times (syndrom bits 8 10)
//  input bit 19 used  2 times (syndrom bits 9 11)
//  input bit 20 used  2 times (syndrom bits 4 6)
//  input bit 21 used  2 times (syndrom bits 5 7)
//  input bit 22 used  2 times (syndrom bits 0 2)
//  input bit 23 used  2 times (syndrom bits 1 3)
//  input bit 24 used  2 times (syndrom bits 0 3)
//  input bit 25 used  2 times (syndrom bits 1 2)
//  input bit 26 used  2 times (syndrom bits 4 7)
//  input bit 27 used  2 times (syndrom bits 5 6)
//  input bit 28 used  2 times (syndrom bits 8 11)
//  input bit 29 used  2 times (syndrom bits 9 10)
//  input bit 30 used  2 times (syndrom bits 12 15)
//  input bit 31 used  2 times (syndrom bits 13 14)
//  input bit 32 used  2 times (syndrom bits 16 19)
//  input bit 33 used  2 times (syndrom bits 17 18)
//  input bit 34 used  2 times (syndrom bits 20 23)
//  input bit 35 used  2 times (syndrom bits 21 22)
//  input bit 36 used  2 times (syndrom bits 17 21)
//  input bit 37 used  2 times (syndrom bits 18 22)
//  input bit 38 used  2 times (syndrom bits 19 23)
//  input bit 39 used  2 times (syndrom bits 16 20)
//  input bit 40 used  2 times (syndrom bits 9 13)
//  input bit 41 used  2 times (syndrom bits 10 14)
//  input bit 42 used  2 times (syndrom bits 11 15)
//  input bit 43 used  2 times (syndrom bits 8 12)
//  input bit 44 used  2 times (syndrom bits 1 5)
//  input bit 45 used  2 times (syndrom bits 2 6)
//  input bit 46 used  2 times (syndrom bits 3 7)
//  input bit 47 used  2 times (syndrom bits 0 4)
function [24-1:0] hamming_code_72_48_f;
    input [48-1:0] in;
    reg [24-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[22]^in[24]^in[47];//4 inputs
        syndrom[ 1] = in[ 0]^in[23]^in[25]^in[44];//4 inputs
        syndrom[ 2] = in[ 1]^in[22]^in[25]^in[45];//4 inputs
        syndrom[ 3] = in[ 1]^in[23]^in[24]^in[46];//4 inputs
        syndrom[ 4] = in[ 2]^in[20]^in[26]^in[47];//4 inputs
        syndrom[ 5] = in[ 2]^in[21]^in[27]^in[44];//4 inputs
        syndrom[ 6] = in[ 3]^in[20]^in[27]^in[45];//4 inputs
        syndrom[ 7] = in[ 3]^in[21]^in[26]^in[46];//4 inputs
        syndrom[ 8] = in[ 4]^in[18]^in[28]^in[43];//4 inputs
        syndrom[ 9] = in[ 4]^in[19]^in[29]^in[40];//4 inputs
        syndrom[10] = in[ 5]^in[18]^in[29]^in[41];//4 inputs
        syndrom[11] = in[ 5]^in[19]^in[28]^in[42];//4 inputs
        syndrom[12] = in[ 6]^in[16]^in[30]^in[43];//4 inputs
        syndrom[13] = in[ 6]^in[17]^in[31]^in[40];//4 inputs
        syndrom[14] = in[ 7]^in[16]^in[31]^in[41];//4 inputs
        syndrom[15] = in[ 7]^in[17]^in[30]^in[42];//4 inputs
        syndrom[16] = in[ 8]^in[14]^in[32]^in[39];//4 inputs
        syndrom[17] = in[ 8]^in[15]^in[33]^in[36];//4 inputs
        syndrom[18] = in[ 9]^in[14]^in[33]^in[37];//4 inputs
        syndrom[19] = in[ 9]^in[15]^in[32]^in[38];//4 inputs
        syndrom[20] = in[10]^in[12]^in[34]^in[39];//4 inputs
        syndrom[21] = in[10]^in[13]^in[35]^in[36];//4 inputs
        syndrom[22] = in[11]^in[12]^in[35]^in[37];//4 inputs
        syndrom[23] = in[11]^in[13]^in[34]^in[38];//4 inputs
        hamming_code_72_48_f = syndrom;
    end
endfunction
wire [24-1:0] stored_data_edc = hamming_code_72_48_f(i_stored_data);
wire [24-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_48_balanced (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [24-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [24-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_72_48_f
//Compute 24 bits Error Detection Code from a 48 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[ 0]: x             x  x             xx             x  (6 inputs)
//  syndrom[ 1]: x              xx              xx              x (6 inputs)
//  syndrom[ 2]: x              x x            x  x            x  (6 inputs)
//  syndrom[ 3]:  x            x x              x x            x  (6 inputs)
//  syndrom[ 4]:  x            x  x            x x              x (6 inputs)
//  syndrom[ 5]:  x             xx             x  x             x (6 inputs)
//  syndrom[ 6]:   x         x      x         x    x         x    (6 inputs)
//  syndrom[ 7]:   x          x    x          x    x          x   (6 inputs)
//  syndrom[ 8]:   x          x     x        x      x        x    (6 inputs)
//  syndrom[ 9]:    x        x     x          x     x        x    (6 inputs)
//  syndrom[10]:    x        x      x        x     x          x   (6 inputs)
//  syndrom[11]:    x         x    x         x      x         x   (6 inputs)
//  syndrom[12]:     x     x          x     x        x     x      (6 inputs)
//  syndrom[13]:     x      x        x      x        x      x     (6 inputs)
//  syndrom[14]:     x      x         x    x          x    x      (6 inputs)
//  syndrom[15]:      x    x         x      x         x    x      (6 inputs)
//  syndrom[16]:      x    x          x    x         x      x     (6 inputs)
//  syndrom[17]:      x     x        x     x          x     x     (6 inputs)
//  syndrom[18]:       x x              x x            x x        (6 inputs)
//  syndrom[19]:       x  x            x  x            x  x       (6 inputs)
//  syndrom[20]:       x  x             xx              xx        (6 inputs)
//  syndrom[21]:        xx             x  x             xx        (6 inputs)
//  syndrom[22]:        xx              xx             x  x       (6 inputs)
//  syndrom[23]:        x x            x x              x x       (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 18 21 22)
//  input bit  9 used  3 times (syndrom bits 19 20 23)
//  input bit 10 used  3 times (syndrom bits 12 15 16)
//  input bit 11 used  3 times (syndrom bits 13 14 17)
//  input bit 12 used  3 times (syndrom bits 6 9 10)
//  input bit 13 used  3 times (syndrom bits 7 8 11)
//  input bit 14 used  3 times (syndrom bits 0 3 4)
//  input bit 15 used  3 times (syndrom bits 1 2 5)
//  input bit 16 used  3 times (syndrom bits 1 3 5)
//  input bit 17 used  3 times (syndrom bits 0 2 4)
//  input bit 18 used  3 times (syndrom bits 7 9 11)
//  input bit 19 used  3 times (syndrom bits 6 8 10)
//  input bit 20 used  3 times (syndrom bits 13 15 17)
//  input bit 21 used  3 times (syndrom bits 12 14 16)
//  input bit 22 used  3 times (syndrom bits 19 21 23)
//  input bit 23 used  3 times (syndrom bits 18 20 22)
//  input bit 24 used  3 times (syndrom bits 20 22 23)
//  input bit 25 used  3 times (syndrom bits 18 19 21)
//  input bit 26 used  3 times (syndrom bits 14 16 17)
//  input bit 27 used  3 times (syndrom bits 12 13 15)
//  input bit 28 used  3 times (syndrom bits 8 10 11)
//  input bit 29 used  3 times (syndrom bits 6 7 9)
//  input bit 30 used  3 times (syndrom bits 2 4 5)
//  input bit 31 used  3 times (syndrom bits 0 1 3)
//  input bit 32 used  3 times (syndrom bits 0 1 4)
//  input bit 33 used  3 times (syndrom bits 2 3 5)
//  input bit 34 used  3 times (syndrom bits 6 7 10)
//  input bit 35 used  3 times (syndrom bits 8 9 11)
//  input bit 36 used  3 times (syndrom bits 12 13 16)
//  input bit 37 used  3 times (syndrom bits 14 15 17)
//  input bit 38 used  3 times (syndrom bits 18 19 22)
//  input bit 39 used  3 times (syndrom bits 20 21 23)
//  input bit 40 used  3 times (syndrom bits 18 20 21)
//  input bit 41 used  3 times (syndrom bits 19 22 23)
//  input bit 42 used  3 times (syndrom bits 12 14 15)
//  input bit 43 used  3 times (syndrom bits 13 16 17)
//  input bit 44 used  3 times (syndrom bits 6 8 9)
//  input bit 45 used  3 times (syndrom bits 7 10 11)
//  input bit 46 used  3 times (syndrom bits 0 2 3)
//  input bit 47 used  3 times (syndrom bits 1 4 5)
function [24-1:0] extended_hamming_code_72_48_f;
    input [48-1:0] in;
    reg [24-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[14]^in[17]^in[31]^in[32]^in[46];//6 inputs
        syndrom[ 1] = in[ 0]^in[15]^in[16]^in[31]^in[32]^in[47];//6 inputs
        syndrom[ 2] = in[ 0]^in[15]^in[17]^in[30]^in[33]^in[46];//6 inputs
        syndrom[ 3] = in[ 1]^in[14]^in[16]^in[31]^in[33]^in[46];//6 inputs
        syndrom[ 4] = in[ 1]^in[14]^in[17]^in[30]^in[32]^in[47];//6 inputs
        syndrom[ 5] = in[ 1]^in[15]^in[16]^in[30]^in[33]^in[47];//6 inputs
        syndrom[ 6] = in[ 2]^in[12]^in[19]^in[29]^in[34]^in[44];//6 inputs
        syndrom[ 7] = in[ 2]^in[13]^in[18]^in[29]^in[34]^in[45];//6 inputs
        syndrom[ 8] = in[ 2]^in[13]^in[19]^in[28]^in[35]^in[44];//6 inputs
        syndrom[ 9] = in[ 3]^in[12]^in[18]^in[29]^in[35]^in[44];//6 inputs
        syndrom[10] = in[ 3]^in[12]^in[19]^in[28]^in[34]^in[45];//6 inputs
        syndrom[11] = in[ 3]^in[13]^in[18]^in[28]^in[35]^in[45];//6 inputs
        syndrom[12] = in[ 4]^in[10]^in[21]^in[27]^in[36]^in[42];//6 inputs
        syndrom[13] = in[ 4]^in[11]^in[20]^in[27]^in[36]^in[43];//6 inputs
        syndrom[14] = in[ 4]^in[11]^in[21]^in[26]^in[37]^in[42];//6 inputs
        syndrom[15] = in[ 5]^in[10]^in[20]^in[27]^in[37]^in[42];//6 inputs
        syndrom[16] = in[ 5]^in[10]^in[21]^in[26]^in[36]^in[43];//6 inputs
        syndrom[17] = in[ 5]^in[11]^in[20]^in[26]^in[37]^in[43];//6 inputs
        syndrom[18] = in[ 6]^in[ 8]^in[23]^in[25]^in[38]^in[40];//6 inputs
        syndrom[19] = in[ 6]^in[ 9]^in[22]^in[25]^in[38]^in[41];//6 inputs
        syndrom[20] = in[ 6]^in[ 9]^in[23]^in[24]^in[39]^in[40];//6 inputs
        syndrom[21] = in[ 7]^in[ 8]^in[22]^in[25]^in[39]^in[40];//6 inputs
        syndrom[22] = in[ 7]^in[ 8]^in[23]^in[24]^in[38]^in[41];//6 inputs
        syndrom[23] = in[ 7]^in[ 9]^in[22]^in[24]^in[39]^in[41];//6 inputs
        extended_hamming_code_72_48_f = syndrom;
    end
endfunction
wire [24-1:0] stored_data_edc = extended_hamming_code_72_48_f(i_stored_data);
wire [24-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_48_balanced (
	input wire [48-1:0] i_write_data, // Data to write to storage
	output reg [24-1:0] o_write_edc, // EDC bits to write to storage
	input wire [48-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [24-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [48-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_72_48_f
//Compute 24 bits Error Detection Code from a 48 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 281474976710656 valid code words out of 4722366482869645213696 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[47]
//  syndrom[ 0]: x             x  x             xx             x  (6 inputs)
//  syndrom[ 1]: x              xx              xx              x (6 inputs)
//  syndrom[ 2]: x              x x            x  x            x  (6 inputs)
//  syndrom[ 3]:  x            x x              x x            x  (6 inputs)
//  syndrom[ 4]:  x            x  x            x x              x (6 inputs)
//  syndrom[ 5]:  x             xx             x  x             x (6 inputs)
//  syndrom[ 6]:   x         x      x         x    x         x    (6 inputs)
//  syndrom[ 7]:   x          x    x          x    x          x   (6 inputs)
//  syndrom[ 8]:   x          x     x        x      x        x    (6 inputs)
//  syndrom[ 9]:    x        x     x          x     x        x    (6 inputs)
//  syndrom[10]:    x        x      x        x     x          x   (6 inputs)
//  syndrom[11]:    x         x    x         x      x         x   (6 inputs)
//  syndrom[12]:     x     x          x     x        x     x      (6 inputs)
//  syndrom[13]:     x      x        x      x        x      x     (6 inputs)
//  syndrom[14]:     x      x         x    x          x    x      (6 inputs)
//  syndrom[15]:      x    x         x      x         x    x      (6 inputs)
//  syndrom[16]:      x    x          x    x         x      x     (6 inputs)
//  syndrom[17]:      x     x        x     x          x     x     (6 inputs)
//  syndrom[18]:       x x              x x            x x        (6 inputs)
//  syndrom[19]:       x  x            x  x            x  x       (6 inputs)
//  syndrom[20]:       x  x             xx              xx        (6 inputs)
//  syndrom[21]:        xx             x  x             xx        (6 inputs)
//  syndrom[22]:        xx              xx             x  x       (6 inputs)
//  syndrom[23]:        x x            x x              x x       (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 18 21 22)
//  input bit  9 used  3 times (syndrom bits 19 20 23)
//  input bit 10 used  3 times (syndrom bits 12 15 16)
//  input bit 11 used  3 times (syndrom bits 13 14 17)
//  input bit 12 used  3 times (syndrom bits 6 9 10)
//  input bit 13 used  3 times (syndrom bits 7 8 11)
//  input bit 14 used  3 times (syndrom bits 0 3 4)
//  input bit 15 used  3 times (syndrom bits 1 2 5)
//  input bit 16 used  3 times (syndrom bits 1 3 5)
//  input bit 17 used  3 times (syndrom bits 0 2 4)
//  input bit 18 used  3 times (syndrom bits 7 9 11)
//  input bit 19 used  3 times (syndrom bits 6 8 10)
//  input bit 20 used  3 times (syndrom bits 13 15 17)
//  input bit 21 used  3 times (syndrom bits 12 14 16)
//  input bit 22 used  3 times (syndrom bits 19 21 23)
//  input bit 23 used  3 times (syndrom bits 18 20 22)
//  input bit 24 used  3 times (syndrom bits 20 22 23)
//  input bit 25 used  3 times (syndrom bits 18 19 21)
//  input bit 26 used  3 times (syndrom bits 14 16 17)
//  input bit 27 used  3 times (syndrom bits 12 13 15)
//  input bit 28 used  3 times (syndrom bits 8 10 11)
//  input bit 29 used  3 times (syndrom bits 6 7 9)
//  input bit 30 used  3 times (syndrom bits 2 4 5)
//  input bit 31 used  3 times (syndrom bits 0 1 3)
//  input bit 32 used  3 times (syndrom bits 0 1 4)
//  input bit 33 used  3 times (syndrom bits 2 3 5)
//  input bit 34 used  3 times (syndrom bits 6 7 10)
//  input bit 35 used  3 times (syndrom bits 8 9 11)
//  input bit 36 used  3 times (syndrom bits 12 13 16)
//  input bit 37 used  3 times (syndrom bits 14 15 17)
//  input bit 38 used  3 times (syndrom bits 18 19 22)
//  input bit 39 used  3 times (syndrom bits 20 21 23)
//  input bit 40 used  3 times (syndrom bits 18 20 21)
//  input bit 41 used  3 times (syndrom bits 19 22 23)
//  input bit 42 used  3 times (syndrom bits 12 14 15)
//  input bit 43 used  3 times (syndrom bits 13 16 17)
//  input bit 44 used  3 times (syndrom bits 6 8 9)
//  input bit 45 used  3 times (syndrom bits 7 10 11)
//  input bit 46 used  3 times (syndrom bits 0 2 3)
//  input bit 47 used  3 times (syndrom bits 1 4 5)
function [24-1:0] extended_hamming_code_72_48_f;
    input [48-1:0] in;
    reg [24-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[14]^in[17]^in[31]^in[32]^in[46];//6 inputs
        syndrom[ 1] = in[ 0]^in[15]^in[16]^in[31]^in[32]^in[47];//6 inputs
        syndrom[ 2] = in[ 0]^in[15]^in[17]^in[30]^in[33]^in[46];//6 inputs
        syndrom[ 3] = in[ 1]^in[14]^in[16]^in[31]^in[33]^in[46];//6 inputs
        syndrom[ 4] = in[ 1]^in[14]^in[17]^in[30]^in[32]^in[47];//6 inputs
        syndrom[ 5] = in[ 1]^in[15]^in[16]^in[30]^in[33]^in[47];//6 inputs
        syndrom[ 6] = in[ 2]^in[12]^in[19]^in[29]^in[34]^in[44];//6 inputs
        syndrom[ 7] = in[ 2]^in[13]^in[18]^in[29]^in[34]^in[45];//6 inputs
        syndrom[ 8] = in[ 2]^in[13]^in[19]^in[28]^in[35]^in[44];//6 inputs
        syndrom[ 9] = in[ 3]^in[12]^in[18]^in[29]^in[35]^in[44];//6 inputs
        syndrom[10] = in[ 3]^in[12]^in[19]^in[28]^in[34]^in[45];//6 inputs
        syndrom[11] = in[ 3]^in[13]^in[18]^in[28]^in[35]^in[45];//6 inputs
        syndrom[12] = in[ 4]^in[10]^in[21]^in[27]^in[36]^in[42];//6 inputs
        syndrom[13] = in[ 4]^in[11]^in[20]^in[27]^in[36]^in[43];//6 inputs
        syndrom[14] = in[ 4]^in[11]^in[21]^in[26]^in[37]^in[42];//6 inputs
        syndrom[15] = in[ 5]^in[10]^in[20]^in[27]^in[37]^in[42];//6 inputs
        syndrom[16] = in[ 5]^in[10]^in[21]^in[26]^in[36]^in[43];//6 inputs
        syndrom[17] = in[ 5]^in[11]^in[20]^in[26]^in[37]^in[43];//6 inputs
        syndrom[18] = in[ 6]^in[ 8]^in[23]^in[25]^in[38]^in[40];//6 inputs
        syndrom[19] = in[ 6]^in[ 9]^in[22]^in[25]^in[38]^in[41];//6 inputs
        syndrom[20] = in[ 6]^in[ 9]^in[23]^in[24]^in[39]^in[40];//6 inputs
        syndrom[21] = in[ 7]^in[ 8]^in[22]^in[25]^in[39]^in[40];//6 inputs
        syndrom[22] = in[ 7]^in[ 8]^in[23]^in[24]^in[38]^in[41];//6 inputs
        syndrom[23] = in[ 7]^in[ 9]^in[22]^in[24]^in[39]^in[41];//6 inputs
        extended_hamming_code_72_48_f = syndrom;
    end
endfunction
function [2+48-1:0] extended_hamming_code_72_48_f_correction_pattern_f;
    input [24-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [48-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {48{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			24'b000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {48{1'b0}};
			end	
			24'b000000000000000000000111: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 0]=1'b1;
			end
			24'b000000000000000000111000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 1]=1'b1;
			end
			24'b000000000000000111000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 2]=1'b1;
			end
			24'b000000000000111000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 3]=1'b1;
			end
			24'b000000000111000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 4]=1'b1;
			end
			24'b000000111000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 5]=1'b1;
			end
			24'b000111000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 6]=1'b1;
			end
			24'b111000000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 7]=1'b1;
			end
			24'b011001000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 8]=1'b1;
			end
			24'b100110000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[ 9]=1'b1;
			end
			24'b000000011001000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[10]=1'b1;
			end
			24'b000000100110000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[11]=1'b1;
			end
			24'b000000000000011001000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[12]=1'b1;
			end
			24'b000000000000100110000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[13]=1'b1;
			end
			24'b000000000000000000011001: begin
				correction_pattern = {48{1'b0}};correction_pattern[14]=1'b1;
			end
			24'b000000000000000000100110: begin
				correction_pattern = {48{1'b0}};correction_pattern[15]=1'b1;
			end
			24'b000000000000000000101010: begin
				correction_pattern = {48{1'b0}};correction_pattern[16]=1'b1;
			end
			24'b000000000000000000010101: begin
				correction_pattern = {48{1'b0}};correction_pattern[17]=1'b1;
			end
			24'b000000000000101010000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[18]=1'b1;
			end
			24'b000000000000010101000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[19]=1'b1;
			end
			24'b000000101010000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[20]=1'b1;
			end
			24'b000000010101000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[21]=1'b1;
			end
			24'b101010000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[22]=1'b1;
			end
			24'b010101000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[23]=1'b1;
			end
			24'b110100000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[24]=1'b1;
			end
			24'b001011000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[25]=1'b1;
			end
			24'b000000110100000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[26]=1'b1;
			end
			24'b000000001011000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[27]=1'b1;
			end
			24'b000000000000110100000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[28]=1'b1;
			end
			24'b000000000000001011000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[29]=1'b1;
			end
			24'b000000000000000000110100: begin
				correction_pattern = {48{1'b0}};correction_pattern[30]=1'b1;
			end
			24'b000000000000000000001011: begin
				correction_pattern = {48{1'b0}};correction_pattern[31]=1'b1;
			end
			24'b000000000000000000010011: begin
				correction_pattern = {48{1'b0}};correction_pattern[32]=1'b1;
			end
			24'b000000000000000000101100: begin
				correction_pattern = {48{1'b0}};correction_pattern[33]=1'b1;
			end
			24'b000000000000010011000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[34]=1'b1;
			end
			24'b000000000000101100000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[35]=1'b1;
			end
			24'b000000010011000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[36]=1'b1;
			end
			24'b000000101100000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[37]=1'b1;
			end
			24'b010011000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[38]=1'b1;
			end
			24'b101100000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[39]=1'b1;
			end
			24'b001101000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[40]=1'b1;
			end
			24'b110010000000000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[41]=1'b1;
			end
			24'b000000001101000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[42]=1'b1;
			end
			24'b000000110010000000000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[43]=1'b1;
			end
			24'b000000000000001101000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[44]=1'b1;
			end
			24'b000000000000110010000000: begin
				correction_pattern = {48{1'b0}};correction_pattern[45]=1'b1;
			end
			24'b000000000000000000001101: begin
				correction_pattern = {48{1'b0}};correction_pattern[46]=1'b1;
			end
			24'b000000000000000000110010: begin
				correction_pattern = {48{1'b0}};correction_pattern[47]=1'b1;
			end
			24'b000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			24'b100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {48{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_72_48_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [24-1:0] stored_data_edc = extended_hamming_code_72_48_f(i_stored_data);
wire [24-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [48-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_72_48_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_64_balanced (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [32-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [32-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_96_64_f
//Compute 32 bits Error Detection Code from a 64 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 79228162514264337593543950336 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[ 0]: x                             x x                              x (4 inputs)
//  syndrom[ 1]: x                              x x                          x    (4 inputs)
//  syndrom[ 2]:  x                            x  x                           x   (4 inputs)
//  syndrom[ 3]:  x                             xx                             x  (4 inputs)
//  syndrom[ 4]:   x                         x     x                            x (4 inputs)
//  syndrom[ 5]:   x                          x     x                        x    (4 inputs)
//  syndrom[ 6]:    x                        x      x                         x   (4 inputs)
//  syndrom[ 7]:    x                         x    x                           x  (4 inputs)
//  syndrom[ 8]:     x                     x         x                      x     (4 inputs)
//  syndrom[ 9]:     x                      x         x                  x        (4 inputs)
//  syndrom[10]:      x                    x          x                   x       (4 inputs)
//  syndrom[11]:      x                     x        x                     x      (4 inputs)
//  syndrom[12]:       x                 x             x                    x     (4 inputs)
//  syndrom[13]:       x                  x             x                x        (4 inputs)
//  syndrom[14]:        x                x              x                 x       (4 inputs)
//  syndrom[15]:        x                 x            x                   x      (4 inputs)
//  syndrom[16]:         x             x                 x              x         (4 inputs)
//  syndrom[17]:         x              x                 x          x            (4 inputs)
//  syndrom[18]:          x            x                  x           x           (4 inputs)
//  syndrom[19]:          x             x                x             x          (4 inputs)
//  syndrom[20]:           x         x                     x            x         (4 inputs)
//  syndrom[21]:           x          x                     x        x            (4 inputs)
//  syndrom[22]:            x        x                      x         x           (4 inputs)
//  syndrom[23]:            x         x                    x           x          (4 inputs)
//  syndrom[24]:             x     x                         x      x             (4 inputs)
//  syndrom[25]:             x      x                         x  x                (4 inputs)
//  syndrom[26]:              x    x                          x   x               (4 inputs)
//  syndrom[27]:              x     x                        x     x              (4 inputs)
//  syndrom[28]:               x x                             x    x             (4 inputs)
//  syndrom[29]:               x  x                             xx                (4 inputs)
//  syndrom[30]:                xx                              x x               (4 inputs)
//  syndrom[31]:                x x                            x   x              (4 inputs)
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 28 30)
//  input bit 17 used  2 times (syndrom bits 29 31)
//  input bit 18 used  2 times (syndrom bits 24 26)
//  input bit 19 used  2 times (syndrom bits 25 27)
//  input bit 20 used  2 times (syndrom bits 20 22)
//  input bit 21 used  2 times (syndrom bits 21 23)
//  input bit 22 used  2 times (syndrom bits 16 18)
//  input bit 23 used  2 times (syndrom bits 17 19)
//  input bit 24 used  2 times (syndrom bits 12 14)
//  input bit 25 used  2 times (syndrom bits 13 15)
//  input bit 26 used  2 times (syndrom bits 8 10)
//  input bit 27 used  2 times (syndrom bits 9 11)
//  input bit 28 used  2 times (syndrom bits 4 6)
//  input bit 29 used  2 times (syndrom bits 5 7)
//  input bit 30 used  2 times (syndrom bits 0 2)
//  input bit 31 used  2 times (syndrom bits 1 3)
//  input bit 32 used  2 times (syndrom bits 0 3)
//  input bit 33 used  2 times (syndrom bits 1 2)
//  input bit 34 used  2 times (syndrom bits 4 7)
//  input bit 35 used  2 times (syndrom bits 5 6)
//  input bit 36 used  2 times (syndrom bits 8 11)
//  input bit 37 used  2 times (syndrom bits 9 10)
//  input bit 38 used  2 times (syndrom bits 12 15)
//  input bit 39 used  2 times (syndrom bits 13 14)
//  input bit 40 used  2 times (syndrom bits 16 19)
//  input bit 41 used  2 times (syndrom bits 17 18)
//  input bit 42 used  2 times (syndrom bits 20 23)
//  input bit 43 used  2 times (syndrom bits 21 22)
//  input bit 44 used  2 times (syndrom bits 24 27)
//  input bit 45 used  2 times (syndrom bits 25 26)
//  input bit 46 used  2 times (syndrom bits 28 31)
//  input bit 47 used  2 times (syndrom bits 29 30)
//  input bit 48 used  2 times (syndrom bits 25 29)
//  input bit 49 used  2 times (syndrom bits 26 30)
//  input bit 50 used  2 times (syndrom bits 27 31)
//  input bit 51 used  2 times (syndrom bits 24 28)
//  input bit 52 used  2 times (syndrom bits 17 21)
//  input bit 53 used  2 times (syndrom bits 18 22)
//  input bit 54 used  2 times (syndrom bits 19 23)
//  input bit 55 used  2 times (syndrom bits 16 20)
//  input bit 56 used  2 times (syndrom bits 9 13)
//  input bit 57 used  2 times (syndrom bits 10 14)
//  input bit 58 used  2 times (syndrom bits 11 15)
//  input bit 59 used  2 times (syndrom bits 8 12)
//  input bit 60 used  2 times (syndrom bits 1 5)
//  input bit 61 used  2 times (syndrom bits 2 6)
//  input bit 62 used  2 times (syndrom bits 3 7)
//  input bit 63 used  2 times (syndrom bits 0 4)
function [32-1:0] hamming_code_96_64_f;
    input [64-1:0] in;
    reg [32-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[30]^in[32]^in[63];//4 inputs
        syndrom[ 1] = in[ 0]^in[31]^in[33]^in[60];//4 inputs
        syndrom[ 2] = in[ 1]^in[30]^in[33]^in[61];//4 inputs
        syndrom[ 3] = in[ 1]^in[31]^in[32]^in[62];//4 inputs
        syndrom[ 4] = in[ 2]^in[28]^in[34]^in[63];//4 inputs
        syndrom[ 5] = in[ 2]^in[29]^in[35]^in[60];//4 inputs
        syndrom[ 6] = in[ 3]^in[28]^in[35]^in[61];//4 inputs
        syndrom[ 7] = in[ 3]^in[29]^in[34]^in[62];//4 inputs
        syndrom[ 8] = in[ 4]^in[26]^in[36]^in[59];//4 inputs
        syndrom[ 9] = in[ 4]^in[27]^in[37]^in[56];//4 inputs
        syndrom[10] = in[ 5]^in[26]^in[37]^in[57];//4 inputs
        syndrom[11] = in[ 5]^in[27]^in[36]^in[58];//4 inputs
        syndrom[12] = in[ 6]^in[24]^in[38]^in[59];//4 inputs
        syndrom[13] = in[ 6]^in[25]^in[39]^in[56];//4 inputs
        syndrom[14] = in[ 7]^in[24]^in[39]^in[57];//4 inputs
        syndrom[15] = in[ 7]^in[25]^in[38]^in[58];//4 inputs
        syndrom[16] = in[ 8]^in[22]^in[40]^in[55];//4 inputs
        syndrom[17] = in[ 8]^in[23]^in[41]^in[52];//4 inputs
        syndrom[18] = in[ 9]^in[22]^in[41]^in[53];//4 inputs
        syndrom[19] = in[ 9]^in[23]^in[40]^in[54];//4 inputs
        syndrom[20] = in[10]^in[20]^in[42]^in[55];//4 inputs
        syndrom[21] = in[10]^in[21]^in[43]^in[52];//4 inputs
        syndrom[22] = in[11]^in[20]^in[43]^in[53];//4 inputs
        syndrom[23] = in[11]^in[21]^in[42]^in[54];//4 inputs
        syndrom[24] = in[12]^in[18]^in[44]^in[51];//4 inputs
        syndrom[25] = in[12]^in[19]^in[45]^in[48];//4 inputs
        syndrom[26] = in[13]^in[18]^in[45]^in[49];//4 inputs
        syndrom[27] = in[13]^in[19]^in[44]^in[50];//4 inputs
        syndrom[28] = in[14]^in[16]^in[46]^in[51];//4 inputs
        syndrom[29] = in[14]^in[17]^in[47]^in[48];//4 inputs
        syndrom[30] = in[15]^in[16]^in[47]^in[49];//4 inputs
        syndrom[31] = in[15]^in[17]^in[46]^in[50];//4 inputs
        hamming_code_96_64_f = syndrom;
    end
endfunction
wire [32-1:0] stored_data_edc = hamming_code_96_64_f(i_stored_data);
wire [32-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_64_balanced (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [32-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [32-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_96_64_f
//Compute 32 bits Error Detection Code from a 64 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 79228162514264337593543950336 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[ 0]: x                   xx                    xx                  x  (6 inputs)
//  syndrom[ 1]: x                   x x                  x  x                x   (6 inputs)
//  syndrom[ 2]: x                    xx                 x    x              x    (6 inputs)
//  syndrom[ 3]:  x                 x   x                x   x                 x  (6 inputs)
//  syndrom[ 4]:  x                 x   x                x   x                 x  (6 inputs)
//  syndrom[ 5]:  x                  xx                    xx                   x (6 inputs)
//  syndrom[ 6]:   x               x     x             x       x             x    (6 inputs)
//  syndrom[ 7]:   x               x     x              x     x               x   (6 inputs)
//  syndrom[ 8]:   x                x  x                  x x                   x (6 inputs)
//  syndrom[ 9]:    x             x       x            x       x             x    (6 inputs)
//  syndrom[10]:    x             x       x            x        x          x      (6 inputs)
//  syndrom[11]:    x              x    x                 xx                    x (6 inputs)
//  syndrom[12]:     x           x         x         x           x         x      (6 inputs)
//  syndrom[13]:     x           x         x          x         x           x     (6 inputs)
//  syndrom[14]:     x            x      x              x      x            x     (6 inputs)
//  syndrom[15]:      x         x           x        x           x         x      (6 inputs)
//  syndrom[16]:      x         x           x        x            x      x        (6 inputs)
//  syndrom[17]:      x          x        x             x     x               x   (6 inputs)
//  syndrom[18]:       x       x             x     x               x     x        (6 inputs)
//  syndrom[19]:       x       x             x      x             x       x       (6 inputs)
//  syndrom[20]:       x        x          x          x          x        x       (6 inputs)
//  syndrom[21]:        x     x               x    x               x     x        (6 inputs)
//  syndrom[22]:        x     x               x    x                x  x          (6 inputs)
//  syndrom[23]:        x      x            x         x         x           x     (6 inputs)
//  syndrom[24]:         x   x                 x x                   xx           (6 inputs)
//  syndrom[25]:         x   x                 x  x                 x   x         (6 inputs)
//  syndrom[26]:         x    x              x      x              x    x         (6 inputs)
//  syndrom[27]:          xx                    x x                 x   x         (6 inputs)
//  syndrom[28]:          x x                   xx                    xx          (6 inputs)
//  syndrom[29]:          x  x                x     x             x       x       (6 inputs)
//  syndrom[30]:           xx                  x  x                  xx           (6 inputs)
//  syndrom[31]:           xx                   xx                   x x          (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 27 30 31)
//  input bit 11 used  3 times (syndrom bits 28 30 31)
//  input bit 12 used  3 times (syndrom bits 24 25 29)
//  input bit 13 used  3 times (syndrom bits 21 22 26)
//  input bit 14 used  3 times (syndrom bits 18 19 23)
//  input bit 15 used  3 times (syndrom bits 15 16 20)
//  input bit 16 used  3 times (syndrom bits 12 13 17)
//  input bit 17 used  3 times (syndrom bits 9 10 14)
//  input bit 18 used  3 times (syndrom bits 6 7 11)
//  input bit 19 used  3 times (syndrom bits 3 4 8)
//  input bit 20 used  3 times (syndrom bits 0 1 5)
//  input bit 21 used  3 times (syndrom bits 0 2 5)
//  input bit 22 used  3 times (syndrom bits 1 2 8)
//  input bit 23 used  3 times (syndrom bits 3 4 11)
//  input bit 24 used  3 times (syndrom bits 6 7 14)
//  input bit 25 used  3 times (syndrom bits 9 10 17)
//  input bit 26 used  3 times (syndrom bits 12 13 20)
//  input bit 27 used  3 times (syndrom bits 15 16 23)
//  input bit 28 used  3 times (syndrom bits 18 19 26)
//  input bit 29 used  3 times (syndrom bits 21 22 29)
//  input bit 30 used  3 times (syndrom bits 24 25 30)
//  input bit 31 used  3 times (syndrom bits 27 28 31)
//  input bit 32 used  3 times (syndrom bits 24 28 31)
//  input bit 33 used  3 times (syndrom bits 25 27 30)
//  input bit 34 used  3 times (syndrom bits 18 21 22)
//  input bit 35 used  3 times (syndrom bits 19 26 29)
//  input bit 36 used  3 times (syndrom bits 12 15 16)
//  input bit 37 used  3 times (syndrom bits 13 20 23)
//  input bit 38 used  3 times (syndrom bits 6 9 10)
//  input bit 39 used  3 times (syndrom bits 7 14 17)
//  input bit 40 used  3 times (syndrom bits 2 3 4)
//  input bit 41 used  3 times (syndrom bits 1 8 11)
//  input bit 42 used  3 times (syndrom bits 0 5 11)
//  input bit 43 used  3 times (syndrom bits 0 5 8)
//  input bit 44 used  3 times (syndrom bits 1 3 4)
//  input bit 45 used  3 times (syndrom bits 2 7 17)
//  input bit 46 used  3 times (syndrom bits 6 9 14)
//  input bit 47 used  3 times (syndrom bits 10 13 23)
//  input bit 48 used  3 times (syndrom bits 12 15 20)
//  input bit 49 used  3 times (syndrom bits 16 19 29)
//  input bit 50 used  3 times (syndrom bits 18 21 26)
//  input bit 51 used  3 times (syndrom bits 22 25 27)
//  input bit 52 used  3 times (syndrom bits 24 30 31)
//  input bit 53 used  3 times (syndrom bits 24 28 30)
//  input bit 54 used  3 times (syndrom bits 22 28 31)
//  input bit 55 used  3 times (syndrom bits 25 26 27)
//  input bit 56 used  3 times (syndrom bits 16 18 21)
//  input bit 57 used  3 times (syndrom bits 19 20 29)
//  input bit 58 used  3 times (syndrom bits 10 12 15)
//  input bit 59 used  3 times (syndrom bits 13 14 23)
//  input bit 60 used  3 times (syndrom bits 2 6 9)
//  input bit 61 used  3 times (syndrom bits 1 7 17)
//  input bit 62 used  3 times (syndrom bits 0 3 4)
//  input bit 63 used  3 times (syndrom bits 5 8 11)
function [32-1:0] extended_hamming_code_96_64_f;
    input [64-1:0] in;
    reg [32-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[20]^in[21]^in[42]^in[43]^in[62];//6 inputs
        syndrom[ 1] = in[ 0]^in[20]^in[22]^in[41]^in[44]^in[61];//6 inputs
        syndrom[ 2] = in[ 0]^in[21]^in[22]^in[40]^in[45]^in[60];//6 inputs
        syndrom[ 3] = in[ 1]^in[19]^in[23]^in[40]^in[44]^in[62];//6 inputs
        syndrom[ 4] = in[ 1]^in[19]^in[23]^in[40]^in[44]^in[62];//6 inputs
        syndrom[ 5] = in[ 1]^in[20]^in[21]^in[42]^in[43]^in[63];//6 inputs
        syndrom[ 6] = in[ 2]^in[18]^in[24]^in[38]^in[46]^in[60];//6 inputs
        syndrom[ 7] = in[ 2]^in[18]^in[24]^in[39]^in[45]^in[61];//6 inputs
        syndrom[ 8] = in[ 2]^in[19]^in[22]^in[41]^in[43]^in[63];//6 inputs
        syndrom[ 9] = in[ 3]^in[17]^in[25]^in[38]^in[46]^in[60];//6 inputs
        syndrom[10] = in[ 3]^in[17]^in[25]^in[38]^in[47]^in[58];//6 inputs
        syndrom[11] = in[ 3]^in[18]^in[23]^in[41]^in[42]^in[63];//6 inputs
        syndrom[12] = in[ 4]^in[16]^in[26]^in[36]^in[48]^in[58];//6 inputs
        syndrom[13] = in[ 4]^in[16]^in[26]^in[37]^in[47]^in[59];//6 inputs
        syndrom[14] = in[ 4]^in[17]^in[24]^in[39]^in[46]^in[59];//6 inputs
        syndrom[15] = in[ 5]^in[15]^in[27]^in[36]^in[48]^in[58];//6 inputs
        syndrom[16] = in[ 5]^in[15]^in[27]^in[36]^in[49]^in[56];//6 inputs
        syndrom[17] = in[ 5]^in[16]^in[25]^in[39]^in[45]^in[61];//6 inputs
        syndrom[18] = in[ 6]^in[14]^in[28]^in[34]^in[50]^in[56];//6 inputs
        syndrom[19] = in[ 6]^in[14]^in[28]^in[35]^in[49]^in[57];//6 inputs
        syndrom[20] = in[ 6]^in[15]^in[26]^in[37]^in[48]^in[57];//6 inputs
        syndrom[21] = in[ 7]^in[13]^in[29]^in[34]^in[50]^in[56];//6 inputs
        syndrom[22] = in[ 7]^in[13]^in[29]^in[34]^in[51]^in[54];//6 inputs
        syndrom[23] = in[ 7]^in[14]^in[27]^in[37]^in[47]^in[59];//6 inputs
        syndrom[24] = in[ 8]^in[12]^in[30]^in[32]^in[52]^in[53];//6 inputs
        syndrom[25] = in[ 8]^in[12]^in[30]^in[33]^in[51]^in[55];//6 inputs
        syndrom[26] = in[ 8]^in[13]^in[28]^in[35]^in[50]^in[55];//6 inputs
        syndrom[27] = in[ 9]^in[10]^in[31]^in[33]^in[51]^in[55];//6 inputs
        syndrom[28] = in[ 9]^in[11]^in[31]^in[32]^in[53]^in[54];//6 inputs
        syndrom[29] = in[ 9]^in[12]^in[29]^in[35]^in[49]^in[57];//6 inputs
        syndrom[30] = in[10]^in[11]^in[30]^in[33]^in[52]^in[53];//6 inputs
        syndrom[31] = in[10]^in[11]^in[31]^in[32]^in[52]^in[54];//6 inputs
        extended_hamming_code_96_64_f = syndrom;
    end
endfunction
wire [32-1:0] stored_data_edc = extended_hamming_code_96_64_f(i_stored_data);
wire [32-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_64_balanced (
	input wire [64-1:0] i_write_data, // Data to write to storage
	output reg [32-1:0] o_write_edc, // EDC bits to write to storage
	input wire [64-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [32-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [64-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_96_64_f
//Compute 32 bits Error Detection Code from a 64 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//There are 18446744073709551616 valid code words out of 79228162514264337593543950336 therefore 99% of errors are detected. 
//Dot graphic view: in[0]...in[63]
//  syndrom[ 0]: x                   xx                    xx                  x  (6 inputs)
//  syndrom[ 1]: x                   x x                  x  x                x   (6 inputs)
//  syndrom[ 2]: x                    xx                 x    x              x    (6 inputs)
//  syndrom[ 3]:  x                 x   x                x   x                 x  (6 inputs)
//  syndrom[ 4]:  x                 x   x                x   x                 x  (6 inputs)
//  syndrom[ 5]:  x                  xx                    xx                   x (6 inputs)
//  syndrom[ 6]:   x               x     x             x       x             x    (6 inputs)
//  syndrom[ 7]:   x               x     x              x     x               x   (6 inputs)
//  syndrom[ 8]:   x                x  x                  x x                   x (6 inputs)
//  syndrom[ 9]:    x             x       x            x       x             x    (6 inputs)
//  syndrom[10]:    x             x       x            x        x          x      (6 inputs)
//  syndrom[11]:    x              x    x                 xx                    x (6 inputs)
//  syndrom[12]:     x           x         x         x           x         x      (6 inputs)
//  syndrom[13]:     x           x         x          x         x           x     (6 inputs)
//  syndrom[14]:     x            x      x              x      x            x     (6 inputs)
//  syndrom[15]:      x         x           x        x           x         x      (6 inputs)
//  syndrom[16]:      x         x           x        x            x      x        (6 inputs)
//  syndrom[17]:      x          x        x             x     x               x   (6 inputs)
//  syndrom[18]:       x       x             x     x               x     x        (6 inputs)
//  syndrom[19]:       x       x             x      x             x       x       (6 inputs)
//  syndrom[20]:       x        x          x          x          x        x       (6 inputs)
//  syndrom[21]:        x     x               x    x               x     x        (6 inputs)
//  syndrom[22]:        x     x               x    x                x  x          (6 inputs)
//  syndrom[23]:        x      x            x         x         x           x     (6 inputs)
//  syndrom[24]:         x   x                 x x                   xx           (6 inputs)
//  syndrom[25]:         x   x                 x  x                 x   x         (6 inputs)
//  syndrom[26]:         x    x              x      x              x    x         (6 inputs)
//  syndrom[27]:          xx                    x x                 x   x         (6 inputs)
//  syndrom[28]:          x x                   xx                    xx          (6 inputs)
//  syndrom[29]:          x  x                x     x             x       x       (6 inputs)
//  syndrom[30]:           xx                  x  x                  xx           (6 inputs)
//  syndrom[31]:           xx                   xx                   x x          (6 inputs)
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 27 30 31)
//  input bit 11 used  3 times (syndrom bits 28 30 31)
//  input bit 12 used  3 times (syndrom bits 24 25 29)
//  input bit 13 used  3 times (syndrom bits 21 22 26)
//  input bit 14 used  3 times (syndrom bits 18 19 23)
//  input bit 15 used  3 times (syndrom bits 15 16 20)
//  input bit 16 used  3 times (syndrom bits 12 13 17)
//  input bit 17 used  3 times (syndrom bits 9 10 14)
//  input bit 18 used  3 times (syndrom bits 6 7 11)
//  input bit 19 used  3 times (syndrom bits 3 4 8)
//  input bit 20 used  3 times (syndrom bits 0 1 5)
//  input bit 21 used  3 times (syndrom bits 0 2 5)
//  input bit 22 used  3 times (syndrom bits 1 2 8)
//  input bit 23 used  3 times (syndrom bits 3 4 11)
//  input bit 24 used  3 times (syndrom bits 6 7 14)
//  input bit 25 used  3 times (syndrom bits 9 10 17)
//  input bit 26 used  3 times (syndrom bits 12 13 20)
//  input bit 27 used  3 times (syndrom bits 15 16 23)
//  input bit 28 used  3 times (syndrom bits 18 19 26)
//  input bit 29 used  3 times (syndrom bits 21 22 29)
//  input bit 30 used  3 times (syndrom bits 24 25 30)
//  input bit 31 used  3 times (syndrom bits 27 28 31)
//  input bit 32 used  3 times (syndrom bits 24 28 31)
//  input bit 33 used  3 times (syndrom bits 25 27 30)
//  input bit 34 used  3 times (syndrom bits 18 21 22)
//  input bit 35 used  3 times (syndrom bits 19 26 29)
//  input bit 36 used  3 times (syndrom bits 12 15 16)
//  input bit 37 used  3 times (syndrom bits 13 20 23)
//  input bit 38 used  3 times (syndrom bits 6 9 10)
//  input bit 39 used  3 times (syndrom bits 7 14 17)
//  input bit 40 used  3 times (syndrom bits 2 3 4)
//  input bit 41 used  3 times (syndrom bits 1 8 11)
//  input bit 42 used  3 times (syndrom bits 0 5 11)
//  input bit 43 used  3 times (syndrom bits 0 5 8)
//  input bit 44 used  3 times (syndrom bits 1 3 4)
//  input bit 45 used  3 times (syndrom bits 2 7 17)
//  input bit 46 used  3 times (syndrom bits 6 9 14)
//  input bit 47 used  3 times (syndrom bits 10 13 23)
//  input bit 48 used  3 times (syndrom bits 12 15 20)
//  input bit 49 used  3 times (syndrom bits 16 19 29)
//  input bit 50 used  3 times (syndrom bits 18 21 26)
//  input bit 51 used  3 times (syndrom bits 22 25 27)
//  input bit 52 used  3 times (syndrom bits 24 30 31)
//  input bit 53 used  3 times (syndrom bits 24 28 30)
//  input bit 54 used  3 times (syndrom bits 22 28 31)
//  input bit 55 used  3 times (syndrom bits 25 26 27)
//  input bit 56 used  3 times (syndrom bits 16 18 21)
//  input bit 57 used  3 times (syndrom bits 19 20 29)
//  input bit 58 used  3 times (syndrom bits 10 12 15)
//  input bit 59 used  3 times (syndrom bits 13 14 23)
//  input bit 60 used  3 times (syndrom bits 2 6 9)
//  input bit 61 used  3 times (syndrom bits 1 7 17)
//  input bit 62 used  3 times (syndrom bits 0 3 4)
//  input bit 63 used  3 times (syndrom bits 5 8 11)
function [32-1:0] extended_hamming_code_96_64_f;
    input [64-1:0] in;
    reg [32-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[20]^in[21]^in[42]^in[43]^in[62];//6 inputs
        syndrom[ 1] = in[ 0]^in[20]^in[22]^in[41]^in[44]^in[61];//6 inputs
        syndrom[ 2] = in[ 0]^in[21]^in[22]^in[40]^in[45]^in[60];//6 inputs
        syndrom[ 3] = in[ 1]^in[19]^in[23]^in[40]^in[44]^in[62];//6 inputs
        syndrom[ 4] = in[ 1]^in[19]^in[23]^in[40]^in[44]^in[62];//6 inputs
        syndrom[ 5] = in[ 1]^in[20]^in[21]^in[42]^in[43]^in[63];//6 inputs
        syndrom[ 6] = in[ 2]^in[18]^in[24]^in[38]^in[46]^in[60];//6 inputs
        syndrom[ 7] = in[ 2]^in[18]^in[24]^in[39]^in[45]^in[61];//6 inputs
        syndrom[ 8] = in[ 2]^in[19]^in[22]^in[41]^in[43]^in[63];//6 inputs
        syndrom[ 9] = in[ 3]^in[17]^in[25]^in[38]^in[46]^in[60];//6 inputs
        syndrom[10] = in[ 3]^in[17]^in[25]^in[38]^in[47]^in[58];//6 inputs
        syndrom[11] = in[ 3]^in[18]^in[23]^in[41]^in[42]^in[63];//6 inputs
        syndrom[12] = in[ 4]^in[16]^in[26]^in[36]^in[48]^in[58];//6 inputs
        syndrom[13] = in[ 4]^in[16]^in[26]^in[37]^in[47]^in[59];//6 inputs
        syndrom[14] = in[ 4]^in[17]^in[24]^in[39]^in[46]^in[59];//6 inputs
        syndrom[15] = in[ 5]^in[15]^in[27]^in[36]^in[48]^in[58];//6 inputs
        syndrom[16] = in[ 5]^in[15]^in[27]^in[36]^in[49]^in[56];//6 inputs
        syndrom[17] = in[ 5]^in[16]^in[25]^in[39]^in[45]^in[61];//6 inputs
        syndrom[18] = in[ 6]^in[14]^in[28]^in[34]^in[50]^in[56];//6 inputs
        syndrom[19] = in[ 6]^in[14]^in[28]^in[35]^in[49]^in[57];//6 inputs
        syndrom[20] = in[ 6]^in[15]^in[26]^in[37]^in[48]^in[57];//6 inputs
        syndrom[21] = in[ 7]^in[13]^in[29]^in[34]^in[50]^in[56];//6 inputs
        syndrom[22] = in[ 7]^in[13]^in[29]^in[34]^in[51]^in[54];//6 inputs
        syndrom[23] = in[ 7]^in[14]^in[27]^in[37]^in[47]^in[59];//6 inputs
        syndrom[24] = in[ 8]^in[12]^in[30]^in[32]^in[52]^in[53];//6 inputs
        syndrom[25] = in[ 8]^in[12]^in[30]^in[33]^in[51]^in[55];//6 inputs
        syndrom[26] = in[ 8]^in[13]^in[28]^in[35]^in[50]^in[55];//6 inputs
        syndrom[27] = in[ 9]^in[10]^in[31]^in[33]^in[51]^in[55];//6 inputs
        syndrom[28] = in[ 9]^in[11]^in[31]^in[32]^in[53]^in[54];//6 inputs
        syndrom[29] = in[ 9]^in[12]^in[29]^in[35]^in[49]^in[57];//6 inputs
        syndrom[30] = in[10]^in[11]^in[30]^in[33]^in[52]^in[53];//6 inputs
        syndrom[31] = in[10]^in[11]^in[31]^in[32]^in[52]^in[54];//6 inputs
        extended_hamming_code_96_64_f = syndrom;
    end
endfunction
function [2+64-1:0] extended_hamming_code_96_64_f_correction_pattern_f;
    input [32-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [64-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {64{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			32'b00000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {64{1'b0}};
			end	
			32'b00000000000000000000000000000111: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 0]=1'b1;
			end
			32'b00000000000000000000000000111000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 1]=1'b1;
			end
			32'b00000000000000000000000111000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 2]=1'b1;
			end
			32'b00000000000000000000111000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 3]=1'b1;
			end
			32'b00000000000000000111000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 4]=1'b1;
			end
			32'b00000000000000111000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 5]=1'b1;
			end
			32'b00000000000111000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 6]=1'b1;
			end
			32'b00000000111000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 7]=1'b1;
			end
			32'b00000111000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 8]=1'b1;
			end
			32'b00111000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[ 9]=1'b1;
			end
			32'b11001000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[10]=1'b1;
			end
			32'b11010000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[11]=1'b1;
			end
			32'b00100011000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[12]=1'b1;
			end
			32'b00000100011000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[13]=1'b1;
			end
			32'b00000000100011000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[14]=1'b1;
			end
			32'b00000000000100011000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[15]=1'b1;
			end
			32'b00000000000000100011000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[16]=1'b1;
			end
			32'b00000000000000000100011000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[17]=1'b1;
			end
			32'b00000000000000000000100011000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[18]=1'b1;
			end
			32'b00000000000000000000000100011000: begin
				correction_pattern = {64{1'b0}};correction_pattern[19]=1'b1;
			end
			32'b00000000000000000000000000100011: begin
				correction_pattern = {64{1'b0}};correction_pattern[20]=1'b1;
			end
			32'b00000000000000000000000000100101: begin
				correction_pattern = {64{1'b0}};correction_pattern[21]=1'b1;
			end
			32'b00000000000000000000000100000110: begin
				correction_pattern = {64{1'b0}};correction_pattern[22]=1'b1;
			end
			32'b00000000000000000000100000011000: begin
				correction_pattern = {64{1'b0}};correction_pattern[23]=1'b1;
			end
			32'b00000000000000000100000011000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[24]=1'b1;
			end
			32'b00000000000000100000011000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[25]=1'b1;
			end
			32'b00000000000100000011000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[26]=1'b1;
			end
			32'b00000000100000011000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[27]=1'b1;
			end
			32'b00000100000011000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[28]=1'b1;
			end
			32'b00100000011000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[29]=1'b1;
			end
			32'b01000011000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[30]=1'b1;
			end
			32'b10011000000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[31]=1'b1;
			end
			32'b10010001000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[32]=1'b1;
			end
			32'b01001010000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[33]=1'b1;
			end
			32'b00000000011001000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[34]=1'b1;
			end
			32'b00100100000010000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[35]=1'b1;
			end
			32'b00000000000000011001000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[36]=1'b1;
			end
			32'b00000000100100000010000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[37]=1'b1;
			end
			32'b00000000000000000000011001000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[38]=1'b1;
			end
			32'b00000000000000100100000010000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[39]=1'b1;
			end
			32'b00000000000000000000000000011100: begin
				correction_pattern = {64{1'b0}};correction_pattern[40]=1'b1;
			end
			32'b00000000000000000000100100000010: begin
				correction_pattern = {64{1'b0}};correction_pattern[41]=1'b1;
			end
			32'b00000000000000000000100000100001: begin
				correction_pattern = {64{1'b0}};correction_pattern[42]=1'b1;
			end
			32'b00000000000000000000000100100001: begin
				correction_pattern = {64{1'b0}};correction_pattern[43]=1'b1;
			end
			32'b00000000000000000000000000011010: begin
				correction_pattern = {64{1'b0}};correction_pattern[44]=1'b1;
			end
			32'b00000000000000100000000010000100: begin
				correction_pattern = {64{1'b0}};correction_pattern[45]=1'b1;
			end
			32'b00000000000000000100001001000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[46]=1'b1;
			end
			32'b00000000100000000010010000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[47]=1'b1;
			end
			32'b00000000000100001001000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[48]=1'b1;
			end
			32'b00100000000010010000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[49]=1'b1;
			end
			32'b00000100001001000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[50]=1'b1;
			end
			32'b00001010010000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[51]=1'b1;
			end
			32'b11000001000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[52]=1'b1;
			end
			32'b01010001000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[53]=1'b1;
			end
			32'b10010000010000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[54]=1'b1;
			end
			32'b00001110000000000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[55]=1'b1;
			end
			32'b00000000001001010000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[56]=1'b1;
			end
			32'b00100000000110000000000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[57]=1'b1;
			end
			32'b00000000000000001001010000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[58]=1'b1;
			end
			32'b00000000100000000110000000000000: begin
				correction_pattern = {64{1'b0}};correction_pattern[59]=1'b1;
			end
			32'b00000000000000000000001001000100: begin
				correction_pattern = {64{1'b0}};correction_pattern[60]=1'b1;
			end
			32'b00000000000000100000000010000010: begin
				correction_pattern = {64{1'b0}};correction_pattern[61]=1'b1;
			end
			32'b00000000000000000000000000011001: begin
				correction_pattern = {64{1'b0}};correction_pattern[62]=1'b1;
			end
			32'b00000000000000000000100100100000: begin
				correction_pattern = {64{1'b0}};correction_pattern[63]=1'b1;
			end
			32'b00000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b00100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b01000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			32'b10000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {64{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_96_64_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [32-1:0] stored_data_edc = extended_hamming_code_96_64_f(i_stored_data);
wire [32-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [64-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_96_64_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_96_balanced (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [48-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [48-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_144_96_f
//Compute 48 bits Error Detection Code from a 96 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used  2 times (syndrom bits 0 1)
//  input bit  1 used  2 times (syndrom bits 2 3)
//  input bit  2 used  2 times (syndrom bits 4 5)
//  input bit  3 used  2 times (syndrom bits 6 7)
//  input bit  4 used  2 times (syndrom bits 8 9)
//  input bit  5 used  2 times (syndrom bits 10 11)
//  input bit  6 used  2 times (syndrom bits 12 13)
//  input bit  7 used  2 times (syndrom bits 14 15)
//  input bit  8 used  2 times (syndrom bits 16 17)
//  input bit  9 used  2 times (syndrom bits 18 19)
//  input bit 10 used  2 times (syndrom bits 20 21)
//  input bit 11 used  2 times (syndrom bits 22 23)
//  input bit 12 used  2 times (syndrom bits 24 25)
//  input bit 13 used  2 times (syndrom bits 26 27)
//  input bit 14 used  2 times (syndrom bits 28 29)
//  input bit 15 used  2 times (syndrom bits 30 31)
//  input bit 16 used  2 times (syndrom bits 32 33)
//  input bit 17 used  2 times (syndrom bits 34 35)
//  input bit 18 used  2 times (syndrom bits 36 37)
//  input bit 19 used  2 times (syndrom bits 38 39)
//  input bit 20 used  2 times (syndrom bits 40 41)
//  input bit 21 used  2 times (syndrom bits 42 43)
//  input bit 22 used  2 times (syndrom bits 44 45)
//  input bit 23 used  2 times (syndrom bits 46 47)
//  input bit 24 used  2 times (syndrom bits 44 46)
//  input bit 25 used  2 times (syndrom bits 45 47)
//  input bit 26 used  2 times (syndrom bits 40 42)
//  input bit 27 used  2 times (syndrom bits 41 43)
//  input bit 28 used  2 times (syndrom bits 36 38)
//  input bit 29 used  2 times (syndrom bits 37 39)
//  input bit 30 used  2 times (syndrom bits 32 34)
//  input bit 31 used  2 times (syndrom bits 33 35)
//  input bit 32 used  2 times (syndrom bits 28 30)
//  input bit 33 used  2 times (syndrom bits 29 31)
//  input bit 34 used  2 times (syndrom bits 24 26)
//  input bit 35 used  2 times (syndrom bits 25 27)
//  input bit 36 used  2 times (syndrom bits 20 22)
//  input bit 37 used  2 times (syndrom bits 21 23)
//  input bit 38 used  2 times (syndrom bits 16 18)
//  input bit 39 used  2 times (syndrom bits 17 19)
//  input bit 40 used  2 times (syndrom bits 12 14)
//  input bit 41 used  2 times (syndrom bits 13 15)
//  input bit 42 used  2 times (syndrom bits 8 10)
//  input bit 43 used  2 times (syndrom bits 9 11)
//  input bit 44 used  2 times (syndrom bits 4 6)
//  input bit 45 used  2 times (syndrom bits 5 7)
//  input bit 46 used  2 times (syndrom bits 0 2)
//  input bit 47 used  2 times (syndrom bits 1 3)
//  input bit 48 used  2 times (syndrom bits 0 3)
//  input bit 49 used  2 times (syndrom bits 1 2)
//  input bit 50 used  2 times (syndrom bits 4 7)
//  input bit 51 used  2 times (syndrom bits 5 6)
//  input bit 52 used  2 times (syndrom bits 8 11)
//  input bit 53 used  2 times (syndrom bits 9 10)
//  input bit 54 used  2 times (syndrom bits 12 15)
//  input bit 55 used  2 times (syndrom bits 13 14)
//  input bit 56 used  2 times (syndrom bits 16 19)
//  input bit 57 used  2 times (syndrom bits 17 18)
//  input bit 58 used  2 times (syndrom bits 20 23)
//  input bit 59 used  2 times (syndrom bits 21 22)
//  input bit 60 used  2 times (syndrom bits 24 27)
//  input bit 61 used  2 times (syndrom bits 25 26)
//  input bit 62 used  2 times (syndrom bits 28 31)
//  input bit 63 used  2 times (syndrom bits 29 30)
//  input bit 64 used  2 times (syndrom bits 32 35)
//  input bit 65 used  2 times (syndrom bits 33 34)
//  input bit 66 used  2 times (syndrom bits 36 39)
//  input bit 67 used  2 times (syndrom bits 37 38)
//  input bit 68 used  2 times (syndrom bits 40 43)
//  input bit 69 used  2 times (syndrom bits 41 42)
//  input bit 70 used  2 times (syndrom bits 44 47)
//  input bit 71 used  2 times (syndrom bits 45 46)
//  input bit 72 used  2 times (syndrom bits 41 45)
//  input bit 73 used  2 times (syndrom bits 42 46)
//  input bit 74 used  2 times (syndrom bits 43 47)
//  input bit 75 used  2 times (syndrom bits 40 44)
//  input bit 76 used  2 times (syndrom bits 33 37)
//  input bit 77 used  2 times (syndrom bits 34 38)
//  input bit 78 used  2 times (syndrom bits 35 39)
//  input bit 79 used  2 times (syndrom bits 32 36)
//  input bit 80 used  2 times (syndrom bits 25 29)
//  input bit 81 used  2 times (syndrom bits 26 30)
//  input bit 82 used  2 times (syndrom bits 27 31)
//  input bit 83 used  2 times (syndrom bits 24 28)
//  input bit 84 used  2 times (syndrom bits 17 21)
//  input bit 85 used  2 times (syndrom bits 18 22)
//  input bit 86 used  2 times (syndrom bits 19 23)
//  input bit 87 used  2 times (syndrom bits 16 20)
//  input bit 88 used  2 times (syndrom bits 9 13)
//  input bit 89 used  2 times (syndrom bits 10 14)
//  input bit 90 used  2 times (syndrom bits 11 15)
//  input bit 91 used  2 times (syndrom bits 8 12)
//  input bit 92 used  2 times (syndrom bits 1 5)
//  input bit 93 used  2 times (syndrom bits 2 6)
//  input bit 94 used  2 times (syndrom bits 3 7)
//  input bit 95 used  2 times (syndrom bits 0 4)
function [48-1:0] hamming_code_144_96_f;
    input [96-1:0] in;
    reg [48-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[46]^in[48]^in[95];//4 inputs
        syndrom[ 1] = in[ 0]^in[47]^in[49]^in[92];//4 inputs
        syndrom[ 2] = in[ 1]^in[46]^in[49]^in[93];//4 inputs
        syndrom[ 3] = in[ 1]^in[47]^in[48]^in[94];//4 inputs
        syndrom[ 4] = in[ 2]^in[44]^in[50]^in[95];//4 inputs
        syndrom[ 5] = in[ 2]^in[45]^in[51]^in[92];//4 inputs
        syndrom[ 6] = in[ 3]^in[44]^in[51]^in[93];//4 inputs
        syndrom[ 7] = in[ 3]^in[45]^in[50]^in[94];//4 inputs
        syndrom[ 8] = in[ 4]^in[42]^in[52]^in[91];//4 inputs
        syndrom[ 9] = in[ 4]^in[43]^in[53]^in[88];//4 inputs
        syndrom[10] = in[ 5]^in[42]^in[53]^in[89];//4 inputs
        syndrom[11] = in[ 5]^in[43]^in[52]^in[90];//4 inputs
        syndrom[12] = in[ 6]^in[40]^in[54]^in[91];//4 inputs
        syndrom[13] = in[ 6]^in[41]^in[55]^in[88];//4 inputs
        syndrom[14] = in[ 7]^in[40]^in[55]^in[89];//4 inputs
        syndrom[15] = in[ 7]^in[41]^in[54]^in[90];//4 inputs
        syndrom[16] = in[ 8]^in[38]^in[56]^in[87];//4 inputs
        syndrom[17] = in[ 8]^in[39]^in[57]^in[84];//4 inputs
        syndrom[18] = in[ 9]^in[38]^in[57]^in[85];//4 inputs
        syndrom[19] = in[ 9]^in[39]^in[56]^in[86];//4 inputs
        syndrom[20] = in[10]^in[36]^in[58]^in[87];//4 inputs
        syndrom[21] = in[10]^in[37]^in[59]^in[84];//4 inputs
        syndrom[22] = in[11]^in[36]^in[59]^in[85];//4 inputs
        syndrom[23] = in[11]^in[37]^in[58]^in[86];//4 inputs
        syndrom[24] = in[12]^in[34]^in[60]^in[83];//4 inputs
        syndrom[25] = in[12]^in[35]^in[61]^in[80];//4 inputs
        syndrom[26] = in[13]^in[34]^in[61]^in[81];//4 inputs
        syndrom[27] = in[13]^in[35]^in[60]^in[82];//4 inputs
        syndrom[28] = in[14]^in[32]^in[62]^in[83];//4 inputs
        syndrom[29] = in[14]^in[33]^in[63]^in[80];//4 inputs
        syndrom[30] = in[15]^in[32]^in[63]^in[81];//4 inputs
        syndrom[31] = in[15]^in[33]^in[62]^in[82];//4 inputs
        syndrom[32] = in[16]^in[30]^in[64]^in[79];//4 inputs
        syndrom[33] = in[16]^in[31]^in[65]^in[76];//4 inputs
        syndrom[34] = in[17]^in[30]^in[65]^in[77];//4 inputs
        syndrom[35] = in[17]^in[31]^in[64]^in[78];//4 inputs
        syndrom[36] = in[18]^in[28]^in[66]^in[79];//4 inputs
        syndrom[37] = in[18]^in[29]^in[67]^in[76];//4 inputs
        syndrom[38] = in[19]^in[28]^in[67]^in[77];//4 inputs
        syndrom[39] = in[19]^in[29]^in[66]^in[78];//4 inputs
        syndrom[40] = in[20]^in[26]^in[68]^in[75];//4 inputs
        syndrom[41] = in[20]^in[27]^in[69]^in[72];//4 inputs
        syndrom[42] = in[21]^in[26]^in[69]^in[73];//4 inputs
        syndrom[43] = in[21]^in[27]^in[68]^in[74];//4 inputs
        syndrom[44] = in[22]^in[24]^in[70]^in[75];//4 inputs
        syndrom[45] = in[22]^in[25]^in[71]^in[72];//4 inputs
        syndrom[46] = in[23]^in[24]^in[71]^in[73];//4 inputs
        syndrom[47] = in[23]^in[25]^in[70]^in[74];//4 inputs
        hamming_code_144_96_f = syndrom;
    end
endfunction
wire [48-1:0] stored_data_edc = hamming_code_144_96_f(i_stored_data);
wire [48-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_96_balanced (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [48-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [48-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_144_96_f
//Compute 48 bits Error Detection Code from a 96 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 42 45 46)
//  input bit 17 used  3 times (syndrom bits 43 44 47)
//  input bit 18 used  3 times (syndrom bits 36 39 40)
//  input bit 19 used  3 times (syndrom bits 37 38 41)
//  input bit 20 used  3 times (syndrom bits 30 33 34)
//  input bit 21 used  3 times (syndrom bits 31 32 35)
//  input bit 22 used  3 times (syndrom bits 24 27 28)
//  input bit 23 used  3 times (syndrom bits 25 26 29)
//  input bit 24 used  3 times (syndrom bits 18 21 22)
//  input bit 25 used  3 times (syndrom bits 19 20 23)
//  input bit 26 used  3 times (syndrom bits 12 15 16)
//  input bit 27 used  3 times (syndrom bits 13 14 17)
//  input bit 28 used  3 times (syndrom bits 6 9 10)
//  input bit 29 used  3 times (syndrom bits 7 8 11)
//  input bit 30 used  3 times (syndrom bits 0 3 4)
//  input bit 31 used  3 times (syndrom bits 1 2 5)
//  input bit 32 used  3 times (syndrom bits 1 3 5)
//  input bit 33 used  3 times (syndrom bits 0 2 4)
//  input bit 34 used  3 times (syndrom bits 7 9 11)
//  input bit 35 used  3 times (syndrom bits 6 8 10)
//  input bit 36 used  3 times (syndrom bits 13 15 17)
//  input bit 37 used  3 times (syndrom bits 12 14 16)
//  input bit 38 used  3 times (syndrom bits 19 21 23)
//  input bit 39 used  3 times (syndrom bits 18 20 22)
//  input bit 40 used  3 times (syndrom bits 25 27 29)
//  input bit 41 used  3 times (syndrom bits 24 26 28)
//  input bit 42 used  3 times (syndrom bits 31 33 35)
//  input bit 43 used  3 times (syndrom bits 30 32 34)
//  input bit 44 used  3 times (syndrom bits 37 39 41)
//  input bit 45 used  3 times (syndrom bits 36 38 40)
//  input bit 46 used  3 times (syndrom bits 43 45 47)
//  input bit 47 used  3 times (syndrom bits 42 44 46)
//  input bit 48 used  3 times (syndrom bits 44 46 47)
//  input bit 49 used  3 times (syndrom bits 42 43 45)
//  input bit 50 used  3 times (syndrom bits 38 40 41)
//  input bit 51 used  3 times (syndrom bits 36 37 39)
//  input bit 52 used  3 times (syndrom bits 32 34 35)
//  input bit 53 used  3 times (syndrom bits 30 31 33)
//  input bit 54 used  3 times (syndrom bits 26 28 29)
//  input bit 55 used  3 times (syndrom bits 24 25 27)
//  input bit 56 used  3 times (syndrom bits 20 22 23)
//  input bit 57 used  3 times (syndrom bits 18 19 21)
//  input bit 58 used  3 times (syndrom bits 14 16 17)
//  input bit 59 used  3 times (syndrom bits 12 13 15)
//  input bit 60 used  3 times (syndrom bits 8 10 11)
//  input bit 61 used  3 times (syndrom bits 6 7 9)
//  input bit 62 used  3 times (syndrom bits 2 4 5)
//  input bit 63 used  3 times (syndrom bits 0 1 3)
//  input bit 64 used  3 times (syndrom bits 0 1 4)
//  input bit 65 used  3 times (syndrom bits 2 3 5)
//  input bit 66 used  3 times (syndrom bits 6 7 10)
//  input bit 67 used  3 times (syndrom bits 8 9 11)
//  input bit 68 used  3 times (syndrom bits 12 13 16)
//  input bit 69 used  3 times (syndrom bits 14 15 17)
//  input bit 70 used  3 times (syndrom bits 18 19 22)
//  input bit 71 used  3 times (syndrom bits 20 21 23)
//  input bit 72 used  3 times (syndrom bits 24 25 28)
//  input bit 73 used  3 times (syndrom bits 26 27 29)
//  input bit 74 used  3 times (syndrom bits 30 31 34)
//  input bit 75 used  3 times (syndrom bits 32 33 35)
//  input bit 76 used  3 times (syndrom bits 36 37 40)
//  input bit 77 used  3 times (syndrom bits 38 39 41)
//  input bit 78 used  3 times (syndrom bits 42 43 46)
//  input bit 79 used  3 times (syndrom bits 44 45 47)
//  input bit 80 used  3 times (syndrom bits 42 44 45)
//  input bit 81 used  3 times (syndrom bits 43 46 47)
//  input bit 82 used  3 times (syndrom bits 36 38 39)
//  input bit 83 used  3 times (syndrom bits 37 40 41)
//  input bit 84 used  3 times (syndrom bits 30 32 33)
//  input bit 85 used  3 times (syndrom bits 31 34 35)
//  input bit 86 used  3 times (syndrom bits 24 26 27)
//  input bit 87 used  3 times (syndrom bits 25 28 29)
//  input bit 88 used  3 times (syndrom bits 18 20 21)
//  input bit 89 used  3 times (syndrom bits 19 22 23)
//  input bit 90 used  3 times (syndrom bits 12 14 15)
//  input bit 91 used  3 times (syndrom bits 13 16 17)
//  input bit 92 used  3 times (syndrom bits 6 8 9)
//  input bit 93 used  3 times (syndrom bits 7 10 11)
//  input bit 94 used  3 times (syndrom bits 0 2 3)
//  input bit 95 used  3 times (syndrom bits 1 4 5)
function [48-1:0] extended_hamming_code_144_96_f;
    input [96-1:0] in;
    reg [48-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[30]^in[33]^in[63]^in[64]^in[94];//6 inputs
        syndrom[ 1] = in[ 0]^in[31]^in[32]^in[63]^in[64]^in[95];//6 inputs
        syndrom[ 2] = in[ 0]^in[31]^in[33]^in[62]^in[65]^in[94];//6 inputs
        syndrom[ 3] = in[ 1]^in[30]^in[32]^in[63]^in[65]^in[94];//6 inputs
        syndrom[ 4] = in[ 1]^in[30]^in[33]^in[62]^in[64]^in[95];//6 inputs
        syndrom[ 5] = in[ 1]^in[31]^in[32]^in[62]^in[65]^in[95];//6 inputs
        syndrom[ 6] = in[ 2]^in[28]^in[35]^in[61]^in[66]^in[92];//6 inputs
        syndrom[ 7] = in[ 2]^in[29]^in[34]^in[61]^in[66]^in[93];//6 inputs
        syndrom[ 8] = in[ 2]^in[29]^in[35]^in[60]^in[67]^in[92];//6 inputs
        syndrom[ 9] = in[ 3]^in[28]^in[34]^in[61]^in[67]^in[92];//6 inputs
        syndrom[10] = in[ 3]^in[28]^in[35]^in[60]^in[66]^in[93];//6 inputs
        syndrom[11] = in[ 3]^in[29]^in[34]^in[60]^in[67]^in[93];//6 inputs
        syndrom[12] = in[ 4]^in[26]^in[37]^in[59]^in[68]^in[90];//6 inputs
        syndrom[13] = in[ 4]^in[27]^in[36]^in[59]^in[68]^in[91];//6 inputs
        syndrom[14] = in[ 4]^in[27]^in[37]^in[58]^in[69]^in[90];//6 inputs
        syndrom[15] = in[ 5]^in[26]^in[36]^in[59]^in[69]^in[90];//6 inputs
        syndrom[16] = in[ 5]^in[26]^in[37]^in[58]^in[68]^in[91];//6 inputs
        syndrom[17] = in[ 5]^in[27]^in[36]^in[58]^in[69]^in[91];//6 inputs
        syndrom[18] = in[ 6]^in[24]^in[39]^in[57]^in[70]^in[88];//6 inputs
        syndrom[19] = in[ 6]^in[25]^in[38]^in[57]^in[70]^in[89];//6 inputs
        syndrom[20] = in[ 6]^in[25]^in[39]^in[56]^in[71]^in[88];//6 inputs
        syndrom[21] = in[ 7]^in[24]^in[38]^in[57]^in[71]^in[88];//6 inputs
        syndrom[22] = in[ 7]^in[24]^in[39]^in[56]^in[70]^in[89];//6 inputs
        syndrom[23] = in[ 7]^in[25]^in[38]^in[56]^in[71]^in[89];//6 inputs
        syndrom[24] = in[ 8]^in[22]^in[41]^in[55]^in[72]^in[86];//6 inputs
        syndrom[25] = in[ 8]^in[23]^in[40]^in[55]^in[72]^in[87];//6 inputs
        syndrom[26] = in[ 8]^in[23]^in[41]^in[54]^in[73]^in[86];//6 inputs
        syndrom[27] = in[ 9]^in[22]^in[40]^in[55]^in[73]^in[86];//6 inputs
        syndrom[28] = in[ 9]^in[22]^in[41]^in[54]^in[72]^in[87];//6 inputs
        syndrom[29] = in[ 9]^in[23]^in[40]^in[54]^in[73]^in[87];//6 inputs
        syndrom[30] = in[10]^in[20]^in[43]^in[53]^in[74]^in[84];//6 inputs
        syndrom[31] = in[10]^in[21]^in[42]^in[53]^in[74]^in[85];//6 inputs
        syndrom[32] = in[10]^in[21]^in[43]^in[52]^in[75]^in[84];//6 inputs
        syndrom[33] = in[11]^in[20]^in[42]^in[53]^in[75]^in[84];//6 inputs
        syndrom[34] = in[11]^in[20]^in[43]^in[52]^in[74]^in[85];//6 inputs
        syndrom[35] = in[11]^in[21]^in[42]^in[52]^in[75]^in[85];//6 inputs
        syndrom[36] = in[12]^in[18]^in[45]^in[51]^in[76]^in[82];//6 inputs
        syndrom[37] = in[12]^in[19]^in[44]^in[51]^in[76]^in[83];//6 inputs
        syndrom[38] = in[12]^in[19]^in[45]^in[50]^in[77]^in[82];//6 inputs
        syndrom[39] = in[13]^in[18]^in[44]^in[51]^in[77]^in[82];//6 inputs
        syndrom[40] = in[13]^in[18]^in[45]^in[50]^in[76]^in[83];//6 inputs
        syndrom[41] = in[13]^in[19]^in[44]^in[50]^in[77]^in[83];//6 inputs
        syndrom[42] = in[14]^in[16]^in[47]^in[49]^in[78]^in[80];//6 inputs
        syndrom[43] = in[14]^in[17]^in[46]^in[49]^in[78]^in[81];//6 inputs
        syndrom[44] = in[14]^in[17]^in[47]^in[48]^in[79]^in[80];//6 inputs
        syndrom[45] = in[15]^in[16]^in[46]^in[49]^in[79]^in[80];//6 inputs
        syndrom[46] = in[15]^in[16]^in[47]^in[48]^in[78]^in[81];//6 inputs
        syndrom[47] = in[15]^in[17]^in[46]^in[48]^in[79]^in[81];//6 inputs
        extended_hamming_code_144_96_f = syndrom;
    end
endfunction
wire [48-1:0] stored_data_edc = extended_hamming_code_144_96_f(i_stored_data);
wire [48-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_96_balanced (
	input wire [96-1:0] i_write_data, // Data to write to storage
	output reg [48-1:0] o_write_edc, // EDC bits to write to storage
	input wire [96-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [48-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [96-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_144_96_f
//Compute 48 bits Error Detection Code from a 96 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit  0 used  3 times (syndrom bits 0 1 2)
//  input bit  1 used  3 times (syndrom bits 3 4 5)
//  input bit  2 used  3 times (syndrom bits 6 7 8)
//  input bit  3 used  3 times (syndrom bits 9 10 11)
//  input bit  4 used  3 times (syndrom bits 12 13 14)
//  input bit  5 used  3 times (syndrom bits 15 16 17)
//  input bit  6 used  3 times (syndrom bits 18 19 20)
//  input bit  7 used  3 times (syndrom bits 21 22 23)
//  input bit  8 used  3 times (syndrom bits 24 25 26)
//  input bit  9 used  3 times (syndrom bits 27 28 29)
//  input bit 10 used  3 times (syndrom bits 30 31 32)
//  input bit 11 used  3 times (syndrom bits 33 34 35)
//  input bit 12 used  3 times (syndrom bits 36 37 38)
//  input bit 13 used  3 times (syndrom bits 39 40 41)
//  input bit 14 used  3 times (syndrom bits 42 43 44)
//  input bit 15 used  3 times (syndrom bits 45 46 47)
//  input bit 16 used  3 times (syndrom bits 42 45 46)
//  input bit 17 used  3 times (syndrom bits 43 44 47)
//  input bit 18 used  3 times (syndrom bits 36 39 40)
//  input bit 19 used  3 times (syndrom bits 37 38 41)
//  input bit 20 used  3 times (syndrom bits 30 33 34)
//  input bit 21 used  3 times (syndrom bits 31 32 35)
//  input bit 22 used  3 times (syndrom bits 24 27 28)
//  input bit 23 used  3 times (syndrom bits 25 26 29)
//  input bit 24 used  3 times (syndrom bits 18 21 22)
//  input bit 25 used  3 times (syndrom bits 19 20 23)
//  input bit 26 used  3 times (syndrom bits 12 15 16)
//  input bit 27 used  3 times (syndrom bits 13 14 17)
//  input bit 28 used  3 times (syndrom bits 6 9 10)
//  input bit 29 used  3 times (syndrom bits 7 8 11)
//  input bit 30 used  3 times (syndrom bits 0 3 4)
//  input bit 31 used  3 times (syndrom bits 1 2 5)
//  input bit 32 used  3 times (syndrom bits 1 3 5)
//  input bit 33 used  3 times (syndrom bits 0 2 4)
//  input bit 34 used  3 times (syndrom bits 7 9 11)
//  input bit 35 used  3 times (syndrom bits 6 8 10)
//  input bit 36 used  3 times (syndrom bits 13 15 17)
//  input bit 37 used  3 times (syndrom bits 12 14 16)
//  input bit 38 used  3 times (syndrom bits 19 21 23)
//  input bit 39 used  3 times (syndrom bits 18 20 22)
//  input bit 40 used  3 times (syndrom bits 25 27 29)
//  input bit 41 used  3 times (syndrom bits 24 26 28)
//  input bit 42 used  3 times (syndrom bits 31 33 35)
//  input bit 43 used  3 times (syndrom bits 30 32 34)
//  input bit 44 used  3 times (syndrom bits 37 39 41)
//  input bit 45 used  3 times (syndrom bits 36 38 40)
//  input bit 46 used  3 times (syndrom bits 43 45 47)
//  input bit 47 used  3 times (syndrom bits 42 44 46)
//  input bit 48 used  3 times (syndrom bits 44 46 47)
//  input bit 49 used  3 times (syndrom bits 42 43 45)
//  input bit 50 used  3 times (syndrom bits 38 40 41)
//  input bit 51 used  3 times (syndrom bits 36 37 39)
//  input bit 52 used  3 times (syndrom bits 32 34 35)
//  input bit 53 used  3 times (syndrom bits 30 31 33)
//  input bit 54 used  3 times (syndrom bits 26 28 29)
//  input bit 55 used  3 times (syndrom bits 24 25 27)
//  input bit 56 used  3 times (syndrom bits 20 22 23)
//  input bit 57 used  3 times (syndrom bits 18 19 21)
//  input bit 58 used  3 times (syndrom bits 14 16 17)
//  input bit 59 used  3 times (syndrom bits 12 13 15)
//  input bit 60 used  3 times (syndrom bits 8 10 11)
//  input bit 61 used  3 times (syndrom bits 6 7 9)
//  input bit 62 used  3 times (syndrom bits 2 4 5)
//  input bit 63 used  3 times (syndrom bits 0 1 3)
//  input bit 64 used  3 times (syndrom bits 0 1 4)
//  input bit 65 used  3 times (syndrom bits 2 3 5)
//  input bit 66 used  3 times (syndrom bits 6 7 10)
//  input bit 67 used  3 times (syndrom bits 8 9 11)
//  input bit 68 used  3 times (syndrom bits 12 13 16)
//  input bit 69 used  3 times (syndrom bits 14 15 17)
//  input bit 70 used  3 times (syndrom bits 18 19 22)
//  input bit 71 used  3 times (syndrom bits 20 21 23)
//  input bit 72 used  3 times (syndrom bits 24 25 28)
//  input bit 73 used  3 times (syndrom bits 26 27 29)
//  input bit 74 used  3 times (syndrom bits 30 31 34)
//  input bit 75 used  3 times (syndrom bits 32 33 35)
//  input bit 76 used  3 times (syndrom bits 36 37 40)
//  input bit 77 used  3 times (syndrom bits 38 39 41)
//  input bit 78 used  3 times (syndrom bits 42 43 46)
//  input bit 79 used  3 times (syndrom bits 44 45 47)
//  input bit 80 used  3 times (syndrom bits 42 44 45)
//  input bit 81 used  3 times (syndrom bits 43 46 47)
//  input bit 82 used  3 times (syndrom bits 36 38 39)
//  input bit 83 used  3 times (syndrom bits 37 40 41)
//  input bit 84 used  3 times (syndrom bits 30 32 33)
//  input bit 85 used  3 times (syndrom bits 31 34 35)
//  input bit 86 used  3 times (syndrom bits 24 26 27)
//  input bit 87 used  3 times (syndrom bits 25 28 29)
//  input bit 88 used  3 times (syndrom bits 18 20 21)
//  input bit 89 used  3 times (syndrom bits 19 22 23)
//  input bit 90 used  3 times (syndrom bits 12 14 15)
//  input bit 91 used  3 times (syndrom bits 13 16 17)
//  input bit 92 used  3 times (syndrom bits 6 8 9)
//  input bit 93 used  3 times (syndrom bits 7 10 11)
//  input bit 94 used  3 times (syndrom bits 0 2 3)
//  input bit 95 used  3 times (syndrom bits 1 4 5)
function [48-1:0] extended_hamming_code_144_96_f;
    input [96-1:0] in;
    reg [48-1:0] syndrom;
    begin
        syndrom[ 0] = in[ 0]^in[30]^in[33]^in[63]^in[64]^in[94];//6 inputs
        syndrom[ 1] = in[ 0]^in[31]^in[32]^in[63]^in[64]^in[95];//6 inputs
        syndrom[ 2] = in[ 0]^in[31]^in[33]^in[62]^in[65]^in[94];//6 inputs
        syndrom[ 3] = in[ 1]^in[30]^in[32]^in[63]^in[65]^in[94];//6 inputs
        syndrom[ 4] = in[ 1]^in[30]^in[33]^in[62]^in[64]^in[95];//6 inputs
        syndrom[ 5] = in[ 1]^in[31]^in[32]^in[62]^in[65]^in[95];//6 inputs
        syndrom[ 6] = in[ 2]^in[28]^in[35]^in[61]^in[66]^in[92];//6 inputs
        syndrom[ 7] = in[ 2]^in[29]^in[34]^in[61]^in[66]^in[93];//6 inputs
        syndrom[ 8] = in[ 2]^in[29]^in[35]^in[60]^in[67]^in[92];//6 inputs
        syndrom[ 9] = in[ 3]^in[28]^in[34]^in[61]^in[67]^in[92];//6 inputs
        syndrom[10] = in[ 3]^in[28]^in[35]^in[60]^in[66]^in[93];//6 inputs
        syndrom[11] = in[ 3]^in[29]^in[34]^in[60]^in[67]^in[93];//6 inputs
        syndrom[12] = in[ 4]^in[26]^in[37]^in[59]^in[68]^in[90];//6 inputs
        syndrom[13] = in[ 4]^in[27]^in[36]^in[59]^in[68]^in[91];//6 inputs
        syndrom[14] = in[ 4]^in[27]^in[37]^in[58]^in[69]^in[90];//6 inputs
        syndrom[15] = in[ 5]^in[26]^in[36]^in[59]^in[69]^in[90];//6 inputs
        syndrom[16] = in[ 5]^in[26]^in[37]^in[58]^in[68]^in[91];//6 inputs
        syndrom[17] = in[ 5]^in[27]^in[36]^in[58]^in[69]^in[91];//6 inputs
        syndrom[18] = in[ 6]^in[24]^in[39]^in[57]^in[70]^in[88];//6 inputs
        syndrom[19] = in[ 6]^in[25]^in[38]^in[57]^in[70]^in[89];//6 inputs
        syndrom[20] = in[ 6]^in[25]^in[39]^in[56]^in[71]^in[88];//6 inputs
        syndrom[21] = in[ 7]^in[24]^in[38]^in[57]^in[71]^in[88];//6 inputs
        syndrom[22] = in[ 7]^in[24]^in[39]^in[56]^in[70]^in[89];//6 inputs
        syndrom[23] = in[ 7]^in[25]^in[38]^in[56]^in[71]^in[89];//6 inputs
        syndrom[24] = in[ 8]^in[22]^in[41]^in[55]^in[72]^in[86];//6 inputs
        syndrom[25] = in[ 8]^in[23]^in[40]^in[55]^in[72]^in[87];//6 inputs
        syndrom[26] = in[ 8]^in[23]^in[41]^in[54]^in[73]^in[86];//6 inputs
        syndrom[27] = in[ 9]^in[22]^in[40]^in[55]^in[73]^in[86];//6 inputs
        syndrom[28] = in[ 9]^in[22]^in[41]^in[54]^in[72]^in[87];//6 inputs
        syndrom[29] = in[ 9]^in[23]^in[40]^in[54]^in[73]^in[87];//6 inputs
        syndrom[30] = in[10]^in[20]^in[43]^in[53]^in[74]^in[84];//6 inputs
        syndrom[31] = in[10]^in[21]^in[42]^in[53]^in[74]^in[85];//6 inputs
        syndrom[32] = in[10]^in[21]^in[43]^in[52]^in[75]^in[84];//6 inputs
        syndrom[33] = in[11]^in[20]^in[42]^in[53]^in[75]^in[84];//6 inputs
        syndrom[34] = in[11]^in[20]^in[43]^in[52]^in[74]^in[85];//6 inputs
        syndrom[35] = in[11]^in[21]^in[42]^in[52]^in[75]^in[85];//6 inputs
        syndrom[36] = in[12]^in[18]^in[45]^in[51]^in[76]^in[82];//6 inputs
        syndrom[37] = in[12]^in[19]^in[44]^in[51]^in[76]^in[83];//6 inputs
        syndrom[38] = in[12]^in[19]^in[45]^in[50]^in[77]^in[82];//6 inputs
        syndrom[39] = in[13]^in[18]^in[44]^in[51]^in[77]^in[82];//6 inputs
        syndrom[40] = in[13]^in[18]^in[45]^in[50]^in[76]^in[83];//6 inputs
        syndrom[41] = in[13]^in[19]^in[44]^in[50]^in[77]^in[83];//6 inputs
        syndrom[42] = in[14]^in[16]^in[47]^in[49]^in[78]^in[80];//6 inputs
        syndrom[43] = in[14]^in[17]^in[46]^in[49]^in[78]^in[81];//6 inputs
        syndrom[44] = in[14]^in[17]^in[47]^in[48]^in[79]^in[80];//6 inputs
        syndrom[45] = in[15]^in[16]^in[46]^in[49]^in[79]^in[80];//6 inputs
        syndrom[46] = in[15]^in[16]^in[47]^in[48]^in[78]^in[81];//6 inputs
        syndrom[47] = in[15]^in[17]^in[46]^in[48]^in[79]^in[81];//6 inputs
        extended_hamming_code_144_96_f = syndrom;
    end
endfunction
function [2+96-1:0] extended_hamming_code_144_96_f_correction_pattern_f;
    input [48-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [96-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {96{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			48'b000000000000000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {96{1'b0}};
			end	
			48'b000000000000000000000000000000000000000000000111: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 0]=1'b1;
			end
			48'b000000000000000000000000000000000000000000111000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 1]=1'b1;
			end
			48'b000000000000000000000000000000000000000111000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 2]=1'b1;
			end
			48'b000000000000000000000000000000000000111000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 3]=1'b1;
			end
			48'b000000000000000000000000000000000111000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 4]=1'b1;
			end
			48'b000000000000000000000000000000111000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 5]=1'b1;
			end
			48'b000000000000000000000000000111000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 6]=1'b1;
			end
			48'b000000000000000000000000111000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 7]=1'b1;
			end
			48'b000000000000000000000111000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 8]=1'b1;
			end
			48'b000000000000000000111000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[ 9]=1'b1;
			end
			48'b000000000000000111000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[10]=1'b1;
			end
			48'b000000000000111000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[11]=1'b1;
			end
			48'b000000000111000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[12]=1'b1;
			end
			48'b000000111000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[13]=1'b1;
			end
			48'b000111000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[14]=1'b1;
			end
			48'b111000000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[15]=1'b1;
			end
			48'b011001000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[16]=1'b1;
			end
			48'b100110000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[17]=1'b1;
			end
			48'b000000011001000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[18]=1'b1;
			end
			48'b000000100110000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[19]=1'b1;
			end
			48'b000000000000011001000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[20]=1'b1;
			end
			48'b000000000000100110000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[21]=1'b1;
			end
			48'b000000000000000000011001000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[22]=1'b1;
			end
			48'b000000000000000000100110000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[23]=1'b1;
			end
			48'b000000000000000000000000011001000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[24]=1'b1;
			end
			48'b000000000000000000000000100110000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[25]=1'b1;
			end
			48'b000000000000000000000000000000011001000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[26]=1'b1;
			end
			48'b000000000000000000000000000000100110000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[27]=1'b1;
			end
			48'b000000000000000000000000000000000000011001000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[28]=1'b1;
			end
			48'b000000000000000000000000000000000000100110000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[29]=1'b1;
			end
			48'b000000000000000000000000000000000000000000011001: begin
				correction_pattern = {96{1'b0}};correction_pattern[30]=1'b1;
			end
			48'b000000000000000000000000000000000000000000100110: begin
				correction_pattern = {96{1'b0}};correction_pattern[31]=1'b1;
			end
			48'b000000000000000000000000000000000000000000101010: begin
				correction_pattern = {96{1'b0}};correction_pattern[32]=1'b1;
			end
			48'b000000000000000000000000000000000000000000010101: begin
				correction_pattern = {96{1'b0}};correction_pattern[33]=1'b1;
			end
			48'b000000000000000000000000000000000000101010000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[34]=1'b1;
			end
			48'b000000000000000000000000000000000000010101000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[35]=1'b1;
			end
			48'b000000000000000000000000000000101010000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[36]=1'b1;
			end
			48'b000000000000000000000000000000010101000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[37]=1'b1;
			end
			48'b000000000000000000000000101010000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[38]=1'b1;
			end
			48'b000000000000000000000000010101000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[39]=1'b1;
			end
			48'b000000000000000000101010000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[40]=1'b1;
			end
			48'b000000000000000000010101000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[41]=1'b1;
			end
			48'b000000000000101010000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[42]=1'b1;
			end
			48'b000000000000010101000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[43]=1'b1;
			end
			48'b000000101010000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[44]=1'b1;
			end
			48'b000000010101000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[45]=1'b1;
			end
			48'b101010000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[46]=1'b1;
			end
			48'b010101000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[47]=1'b1;
			end
			48'b110100000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[48]=1'b1;
			end
			48'b001011000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[49]=1'b1;
			end
			48'b000000110100000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[50]=1'b1;
			end
			48'b000000001011000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[51]=1'b1;
			end
			48'b000000000000110100000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[52]=1'b1;
			end
			48'b000000000000001011000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[53]=1'b1;
			end
			48'b000000000000000000110100000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[54]=1'b1;
			end
			48'b000000000000000000001011000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[55]=1'b1;
			end
			48'b000000000000000000000000110100000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[56]=1'b1;
			end
			48'b000000000000000000000000001011000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[57]=1'b1;
			end
			48'b000000000000000000000000000000110100000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[58]=1'b1;
			end
			48'b000000000000000000000000000000001011000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[59]=1'b1;
			end
			48'b000000000000000000000000000000000000110100000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[60]=1'b1;
			end
			48'b000000000000000000000000000000000000001011000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[61]=1'b1;
			end
			48'b000000000000000000000000000000000000000000110100: begin
				correction_pattern = {96{1'b0}};correction_pattern[62]=1'b1;
			end
			48'b000000000000000000000000000000000000000000001011: begin
				correction_pattern = {96{1'b0}};correction_pattern[63]=1'b1;
			end
			48'b000000000000000000000000000000000000000000010011: begin
				correction_pattern = {96{1'b0}};correction_pattern[64]=1'b1;
			end
			48'b000000000000000000000000000000000000000000101100: begin
				correction_pattern = {96{1'b0}};correction_pattern[65]=1'b1;
			end
			48'b000000000000000000000000000000000000010011000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[66]=1'b1;
			end
			48'b000000000000000000000000000000000000101100000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[67]=1'b1;
			end
			48'b000000000000000000000000000000010011000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[68]=1'b1;
			end
			48'b000000000000000000000000000000101100000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[69]=1'b1;
			end
			48'b000000000000000000000000010011000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[70]=1'b1;
			end
			48'b000000000000000000000000101100000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[71]=1'b1;
			end
			48'b000000000000000000010011000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[72]=1'b1;
			end
			48'b000000000000000000101100000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[73]=1'b1;
			end
			48'b000000000000010011000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[74]=1'b1;
			end
			48'b000000000000101100000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[75]=1'b1;
			end
			48'b000000010011000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[76]=1'b1;
			end
			48'b000000101100000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[77]=1'b1;
			end
			48'b010011000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[78]=1'b1;
			end
			48'b101100000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[79]=1'b1;
			end
			48'b001101000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[80]=1'b1;
			end
			48'b110010000000000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[81]=1'b1;
			end
			48'b000000001101000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[82]=1'b1;
			end
			48'b000000110010000000000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[83]=1'b1;
			end
			48'b000000000000001101000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[84]=1'b1;
			end
			48'b000000000000110010000000000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[85]=1'b1;
			end
			48'b000000000000000000001101000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[86]=1'b1;
			end
			48'b000000000000000000110010000000000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[87]=1'b1;
			end
			48'b000000000000000000000000001101000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[88]=1'b1;
			end
			48'b000000000000000000000000110010000000000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[89]=1'b1;
			end
			48'b000000000000000000000000000000001101000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[90]=1'b1;
			end
			48'b000000000000000000000000000000110010000000000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[91]=1'b1;
			end
			48'b000000000000000000000000000000000000001101000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[92]=1'b1;
			end
			48'b000000000000000000000000000000000000110010000000: begin
				correction_pattern = {96{1'b0}};correction_pattern[93]=1'b1;
			end
			48'b000000000000000000000000000000000000000000001101: begin
				correction_pattern = {96{1'b0}};correction_pattern[94]=1'b1;
			end
			48'b000000000000000000000000000000000000000000110010: begin
				correction_pattern = {96{1'b0}};correction_pattern[95]=1'b1;
			end
			48'b000000000000000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000000100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000001000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000010000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000000100000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000001000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000010000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000000100000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000001000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000010000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b000100000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b001000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b010000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			48'b100000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {96{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_144_96_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [48-1:0] stored_data_edc = extended_hamming_code_144_96_f(i_stored_data);
wire [48-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [96-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_144_96_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule

module edc_hc_128_balanced (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [64-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [64-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//hamming_code_192_128_f
//Compute 64 bits Error Detection Code from a 128 bits input.
//The EDC is a hamming code capable of detecting any 1 and 2 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used  2 times (syndrom bits 0 1)
//  input bit   1 used  2 times (syndrom bits 2 3)
//  input bit   2 used  2 times (syndrom bits 4 5)
//  input bit   3 used  2 times (syndrom bits 6 7)
//  input bit   4 used  2 times (syndrom bits 8 9)
//  input bit   5 used  2 times (syndrom bits 10 11)
//  input bit   6 used  2 times (syndrom bits 12 13)
//  input bit   7 used  2 times (syndrom bits 14 15)
//  input bit   8 used  2 times (syndrom bits 16 17)
//  input bit   9 used  2 times (syndrom bits 18 19)
//  input bit  10 used  2 times (syndrom bits 20 21)
//  input bit  11 used  2 times (syndrom bits 22 23)
//  input bit  12 used  2 times (syndrom bits 24 25)
//  input bit  13 used  2 times (syndrom bits 26 27)
//  input bit  14 used  2 times (syndrom bits 28 29)
//  input bit  15 used  2 times (syndrom bits 30 31)
//  input bit  16 used  2 times (syndrom bits 32 33)
//  input bit  17 used  2 times (syndrom bits 34 35)
//  input bit  18 used  2 times (syndrom bits 36 37)
//  input bit  19 used  2 times (syndrom bits 38 39)
//  input bit  20 used  2 times (syndrom bits 40 41)
//  input bit  21 used  2 times (syndrom bits 42 43)
//  input bit  22 used  2 times (syndrom bits 44 45)
//  input bit  23 used  2 times (syndrom bits 46 47)
//  input bit  24 used  2 times (syndrom bits 48 49)
//  input bit  25 used  2 times (syndrom bits 50 51)
//  input bit  26 used  2 times (syndrom bits 52 53)
//  input bit  27 used  2 times (syndrom bits 54 55)
//  input bit  28 used  2 times (syndrom bits 56 57)
//  input bit  29 used  2 times (syndrom bits 58 59)
//  input bit  30 used  2 times (syndrom bits 60 61)
//  input bit  31 used  2 times (syndrom bits 62 63)
//  input bit  32 used  2 times (syndrom bits 60 62)
//  input bit  33 used  2 times (syndrom bits 61 63)
//  input bit  34 used  2 times (syndrom bits 56 58)
//  input bit  35 used  2 times (syndrom bits 57 59)
//  input bit  36 used  2 times (syndrom bits 52 54)
//  input bit  37 used  2 times (syndrom bits 53 55)
//  input bit  38 used  2 times (syndrom bits 48 50)
//  input bit  39 used  2 times (syndrom bits 49 51)
//  input bit  40 used  2 times (syndrom bits 44 46)
//  input bit  41 used  2 times (syndrom bits 45 47)
//  input bit  42 used  2 times (syndrom bits 40 42)
//  input bit  43 used  2 times (syndrom bits 41 43)
//  input bit  44 used  2 times (syndrom bits 36 38)
//  input bit  45 used  2 times (syndrom bits 37 39)
//  input bit  46 used  2 times (syndrom bits 32 34)
//  input bit  47 used  2 times (syndrom bits 33 35)
//  input bit  48 used  2 times (syndrom bits 28 30)
//  input bit  49 used  2 times (syndrom bits 29 31)
//  input bit  50 used  2 times (syndrom bits 24 26)
//  input bit  51 used  2 times (syndrom bits 25 27)
//  input bit  52 used  2 times (syndrom bits 20 22)
//  input bit  53 used  2 times (syndrom bits 21 23)
//  input bit  54 used  2 times (syndrom bits 16 18)
//  input bit  55 used  2 times (syndrom bits 17 19)
//  input bit  56 used  2 times (syndrom bits 12 14)
//  input bit  57 used  2 times (syndrom bits 13 15)
//  input bit  58 used  2 times (syndrom bits 8 10)
//  input bit  59 used  2 times (syndrom bits 9 11)
//  input bit  60 used  2 times (syndrom bits 4 6)
//  input bit  61 used  2 times (syndrom bits 5 7)
//  input bit  62 used  2 times (syndrom bits 0 2)
//  input bit  63 used  2 times (syndrom bits 1 3)
//  input bit  64 used  2 times (syndrom bits 0 3)
//  input bit  65 used  2 times (syndrom bits 1 2)
//  input bit  66 used  2 times (syndrom bits 4 7)
//  input bit  67 used  2 times (syndrom bits 5 6)
//  input bit  68 used  2 times (syndrom bits 8 11)
//  input bit  69 used  2 times (syndrom bits 9 10)
//  input bit  70 used  2 times (syndrom bits 12 15)
//  input bit  71 used  2 times (syndrom bits 13 14)
//  input bit  72 used  2 times (syndrom bits 16 19)
//  input bit  73 used  2 times (syndrom bits 17 18)
//  input bit  74 used  2 times (syndrom bits 20 23)
//  input bit  75 used  2 times (syndrom bits 21 22)
//  input bit  76 used  2 times (syndrom bits 24 27)
//  input bit  77 used  2 times (syndrom bits 25 26)
//  input bit  78 used  2 times (syndrom bits 28 31)
//  input bit  79 used  2 times (syndrom bits 29 30)
//  input bit  80 used  2 times (syndrom bits 32 35)
//  input bit  81 used  2 times (syndrom bits 33 34)
//  input bit  82 used  2 times (syndrom bits 36 39)
//  input bit  83 used  2 times (syndrom bits 37 38)
//  input bit  84 used  2 times (syndrom bits 40 43)
//  input bit  85 used  2 times (syndrom bits 41 42)
//  input bit  86 used  2 times (syndrom bits 44 47)
//  input bit  87 used  2 times (syndrom bits 45 46)
//  input bit  88 used  2 times (syndrom bits 48 51)
//  input bit  89 used  2 times (syndrom bits 49 50)
//  input bit  90 used  2 times (syndrom bits 52 55)
//  input bit  91 used  2 times (syndrom bits 53 54)
//  input bit  92 used  2 times (syndrom bits 56 59)
//  input bit  93 used  2 times (syndrom bits 57 58)
//  input bit  94 used  2 times (syndrom bits 60 63)
//  input bit  95 used  2 times (syndrom bits 61 62)
//  input bit  96 used  2 times (syndrom bits 57 61)
//  input bit  97 used  2 times (syndrom bits 58 62)
//  input bit  98 used  2 times (syndrom bits 59 63)
//  input bit  99 used  2 times (syndrom bits 56 60)
//  input bit 100 used  2 times (syndrom bits 49 53)
//  input bit 101 used  2 times (syndrom bits 50 54)
//  input bit 102 used  2 times (syndrom bits 51 55)
//  input bit 103 used  2 times (syndrom bits 48 52)
//  input bit 104 used  2 times (syndrom bits 41 45)
//  input bit 105 used  2 times (syndrom bits 42 46)
//  input bit 106 used  2 times (syndrom bits 43 47)
//  input bit 107 used  2 times (syndrom bits 40 44)
//  input bit 108 used  2 times (syndrom bits 33 37)
//  input bit 109 used  2 times (syndrom bits 34 38)
//  input bit 110 used  2 times (syndrom bits 35 39)
//  input bit 111 used  2 times (syndrom bits 32 36)
//  input bit 112 used  2 times (syndrom bits 25 29)
//  input bit 113 used  2 times (syndrom bits 26 30)
//  input bit 114 used  2 times (syndrom bits 27 31)
//  input bit 115 used  2 times (syndrom bits 24 28)
//  input bit 116 used  2 times (syndrom bits 17 21)
//  input bit 117 used  2 times (syndrom bits 18 22)
//  input bit 118 used  2 times (syndrom bits 19 23)
//  input bit 119 used  2 times (syndrom bits 16 20)
//  input bit 120 used  2 times (syndrom bits 9 13)
//  input bit 121 used  2 times (syndrom bits 10 14)
//  input bit 122 used  2 times (syndrom bits 11 15)
//  input bit 123 used  2 times (syndrom bits 8 12)
//  input bit 124 used  2 times (syndrom bits 1 5)
//  input bit 125 used  2 times (syndrom bits 2 6)
//  input bit 126 used  2 times (syndrom bits 3 7)
//  input bit 127 used  2 times (syndrom bits 0 4)
function [64-1:0] hamming_code_192_128_f;
    input [128-1:0] in;
    reg [64-1:0] syndrom;
    begin
        syndrom[ 0] = in[  0]^in[ 62]^in[ 64]^in[127];//4 inputs
        syndrom[ 1] = in[  0]^in[ 63]^in[ 65]^in[124];//4 inputs
        syndrom[ 2] = in[  1]^in[ 62]^in[ 65]^in[125];//4 inputs
        syndrom[ 3] = in[  1]^in[ 63]^in[ 64]^in[126];//4 inputs
        syndrom[ 4] = in[  2]^in[ 60]^in[ 66]^in[127];//4 inputs
        syndrom[ 5] = in[  2]^in[ 61]^in[ 67]^in[124];//4 inputs
        syndrom[ 6] = in[  3]^in[ 60]^in[ 67]^in[125];//4 inputs
        syndrom[ 7] = in[  3]^in[ 61]^in[ 66]^in[126];//4 inputs
        syndrom[ 8] = in[  4]^in[ 58]^in[ 68]^in[123];//4 inputs
        syndrom[ 9] = in[  4]^in[ 59]^in[ 69]^in[120];//4 inputs
        syndrom[10] = in[  5]^in[ 58]^in[ 69]^in[121];//4 inputs
        syndrom[11] = in[  5]^in[ 59]^in[ 68]^in[122];//4 inputs
        syndrom[12] = in[  6]^in[ 56]^in[ 70]^in[123];//4 inputs
        syndrom[13] = in[  6]^in[ 57]^in[ 71]^in[120];//4 inputs
        syndrom[14] = in[  7]^in[ 56]^in[ 71]^in[121];//4 inputs
        syndrom[15] = in[  7]^in[ 57]^in[ 70]^in[122];//4 inputs
        syndrom[16] = in[  8]^in[ 54]^in[ 72]^in[119];//4 inputs
        syndrom[17] = in[  8]^in[ 55]^in[ 73]^in[116];//4 inputs
        syndrom[18] = in[  9]^in[ 54]^in[ 73]^in[117];//4 inputs
        syndrom[19] = in[  9]^in[ 55]^in[ 72]^in[118];//4 inputs
        syndrom[20] = in[ 10]^in[ 52]^in[ 74]^in[119];//4 inputs
        syndrom[21] = in[ 10]^in[ 53]^in[ 75]^in[116];//4 inputs
        syndrom[22] = in[ 11]^in[ 52]^in[ 75]^in[117];//4 inputs
        syndrom[23] = in[ 11]^in[ 53]^in[ 74]^in[118];//4 inputs
        syndrom[24] = in[ 12]^in[ 50]^in[ 76]^in[115];//4 inputs
        syndrom[25] = in[ 12]^in[ 51]^in[ 77]^in[112];//4 inputs
        syndrom[26] = in[ 13]^in[ 50]^in[ 77]^in[113];//4 inputs
        syndrom[27] = in[ 13]^in[ 51]^in[ 76]^in[114];//4 inputs
        syndrom[28] = in[ 14]^in[ 48]^in[ 78]^in[115];//4 inputs
        syndrom[29] = in[ 14]^in[ 49]^in[ 79]^in[112];//4 inputs
        syndrom[30] = in[ 15]^in[ 48]^in[ 79]^in[113];//4 inputs
        syndrom[31] = in[ 15]^in[ 49]^in[ 78]^in[114];//4 inputs
        syndrom[32] = in[ 16]^in[ 46]^in[ 80]^in[111];//4 inputs
        syndrom[33] = in[ 16]^in[ 47]^in[ 81]^in[108];//4 inputs
        syndrom[34] = in[ 17]^in[ 46]^in[ 81]^in[109];//4 inputs
        syndrom[35] = in[ 17]^in[ 47]^in[ 80]^in[110];//4 inputs
        syndrom[36] = in[ 18]^in[ 44]^in[ 82]^in[111];//4 inputs
        syndrom[37] = in[ 18]^in[ 45]^in[ 83]^in[108];//4 inputs
        syndrom[38] = in[ 19]^in[ 44]^in[ 83]^in[109];//4 inputs
        syndrom[39] = in[ 19]^in[ 45]^in[ 82]^in[110];//4 inputs
        syndrom[40] = in[ 20]^in[ 42]^in[ 84]^in[107];//4 inputs
        syndrom[41] = in[ 20]^in[ 43]^in[ 85]^in[104];//4 inputs
        syndrom[42] = in[ 21]^in[ 42]^in[ 85]^in[105];//4 inputs
        syndrom[43] = in[ 21]^in[ 43]^in[ 84]^in[106];//4 inputs
        syndrom[44] = in[ 22]^in[ 40]^in[ 86]^in[107];//4 inputs
        syndrom[45] = in[ 22]^in[ 41]^in[ 87]^in[104];//4 inputs
        syndrom[46] = in[ 23]^in[ 40]^in[ 87]^in[105];//4 inputs
        syndrom[47] = in[ 23]^in[ 41]^in[ 86]^in[106];//4 inputs
        syndrom[48] = in[ 24]^in[ 38]^in[ 88]^in[103];//4 inputs
        syndrom[49] = in[ 24]^in[ 39]^in[ 89]^in[100];//4 inputs
        syndrom[50] = in[ 25]^in[ 38]^in[ 89]^in[101];//4 inputs
        syndrom[51] = in[ 25]^in[ 39]^in[ 88]^in[102];//4 inputs
        syndrom[52] = in[ 26]^in[ 36]^in[ 90]^in[103];//4 inputs
        syndrom[53] = in[ 26]^in[ 37]^in[ 91]^in[100];//4 inputs
        syndrom[54] = in[ 27]^in[ 36]^in[ 91]^in[101];//4 inputs
        syndrom[55] = in[ 27]^in[ 37]^in[ 90]^in[102];//4 inputs
        syndrom[56] = in[ 28]^in[ 34]^in[ 92]^in[ 99];//4 inputs
        syndrom[57] = in[ 28]^in[ 35]^in[ 93]^in[ 96];//4 inputs
        syndrom[58] = in[ 29]^in[ 34]^in[ 93]^in[ 97];//4 inputs
        syndrom[59] = in[ 29]^in[ 35]^in[ 92]^in[ 98];//4 inputs
        syndrom[60] = in[ 30]^in[ 32]^in[ 94]^in[ 99];//4 inputs
        syndrom[61] = in[ 30]^in[ 33]^in[ 95]^in[ 96];//4 inputs
        syndrom[62] = in[ 31]^in[ 32]^in[ 95]^in[ 97];//4 inputs
        syndrom[63] = in[ 31]^in[ 33]^in[ 94]^in[ 98];//4 inputs
        hamming_code_192_128_f = syndrom;
    end
endfunction
wire [64-1:0] stored_data_edc = hamming_code_192_128_f(i_stored_data);
wire [64-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module edc_ehc_128_balanced (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [64-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [64-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg o_detection //indication that an error is detected
);
//extended_hamming_code_192_128_f
//Compute 64 bits Error Detection Code from a 128 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used  3 times (syndrom bits 0 1 2)
//  input bit   1 used  3 times (syndrom bits 3 4 5)
//  input bit   2 used  3 times (syndrom bits 6 7 8)
//  input bit   3 used  3 times (syndrom bits 9 10 11)
//  input bit   4 used  3 times (syndrom bits 12 13 14)
//  input bit   5 used  3 times (syndrom bits 15 16 17)
//  input bit   6 used  3 times (syndrom bits 18 19 20)
//  input bit   7 used  3 times (syndrom bits 21 22 23)
//  input bit   8 used  3 times (syndrom bits 24 25 26)
//  input bit   9 used  3 times (syndrom bits 27 28 29)
//  input bit  10 used  3 times (syndrom bits 30 31 32)
//  input bit  11 used  3 times (syndrom bits 33 34 35)
//  input bit  12 used  3 times (syndrom bits 36 37 38)
//  input bit  13 used  3 times (syndrom bits 39 40 41)
//  input bit  14 used  3 times (syndrom bits 42 43 44)
//  input bit  15 used  3 times (syndrom bits 45 46 47)
//  input bit  16 used  3 times (syndrom bits 48 49 50)
//  input bit  17 used  3 times (syndrom bits 51 52 53)
//  input bit  18 used  3 times (syndrom bits 54 55 56)
//  input bit  19 used  3 times (syndrom bits 57 58 59)
//  input bit  20 used  3 times (syndrom bits 60 61 62)
//  input bit  21 used  3 times (syndrom bits 60 61 63)
//  input bit  22 used  3 times (syndrom bits 57 62 63)
//  input bit  23 used  3 times (syndrom bits 54 58 59)
//  input bit  24 used  3 times (syndrom bits 51 55 56)
//  input bit  25 used  3 times (syndrom bits 48 52 53)
//  input bit  26 used  3 times (syndrom bits 45 49 50)
//  input bit  27 used  3 times (syndrom bits 42 46 47)
//  input bit  28 used  3 times (syndrom bits 39 43 44)
//  input bit  29 used  3 times (syndrom bits 36 40 41)
//  input bit  30 used  3 times (syndrom bits 33 37 38)
//  input bit  31 used  3 times (syndrom bits 30 34 35)
//  input bit  32 used  3 times (syndrom bits 27 31 32)
//  input bit  33 used  3 times (syndrom bits 24 28 29)
//  input bit  34 used  3 times (syndrom bits 21 25 26)
//  input bit  35 used  3 times (syndrom bits 18 22 23)
//  input bit  36 used  3 times (syndrom bits 15 19 20)
//  input bit  37 used  3 times (syndrom bits 12 16 17)
//  input bit  38 used  3 times (syndrom bits 9 13 14)
//  input bit  39 used  3 times (syndrom bits 6 10 11)
//  input bit  40 used  3 times (syndrom bits 3 7 8)
//  input bit  41 used  3 times (syndrom bits 0 4 5)
//  input bit  42 used  3 times (syndrom bits 1 2 4)
//  input bit  43 used  3 times (syndrom bits 1 2 5)
//  input bit  44 used  3 times (syndrom bits 0 7 8)
//  input bit  45 used  3 times (syndrom bits 3 10 11)
//  input bit  46 used  3 times (syndrom bits 6 13 14)
//  input bit  47 used  3 times (syndrom bits 9 16 17)
//  input bit  48 used  3 times (syndrom bits 12 19 20)
//  input bit  49 used  3 times (syndrom bits 15 22 23)
//  input bit  50 used  3 times (syndrom bits 18 25 26)
//  input bit  51 used  3 times (syndrom bits 21 28 29)
//  input bit  52 used  3 times (syndrom bits 24 31 32)
//  input bit  53 used  3 times (syndrom bits 27 34 35)
//  input bit  54 used  3 times (syndrom bits 30 37 38)
//  input bit  55 used  3 times (syndrom bits 33 40 41)
//  input bit  56 used  3 times (syndrom bits 36 43 44)
//  input bit  57 used  3 times (syndrom bits 39 46 47)
//  input bit  58 used  3 times (syndrom bits 42 49 50)
//  input bit  59 used  3 times (syndrom bits 45 52 53)
//  input bit  60 used  3 times (syndrom bits 48 55 56)
//  input bit  61 used  3 times (syndrom bits 51 58 59)
//  input bit  62 used  3 times (syndrom bits 54 62 63)
//  input bit  63 used  3 times (syndrom bits 57 60 61)
//  input bit  64 used  3 times (syndrom bits 54 57 60)
//  input bit  65 used  3 times (syndrom bits 61 62 63)
//  input bit  66 used  3 times (syndrom bits 48 51 58)
//  input bit  67 used  3 times (syndrom bits 55 56 59)
//  input bit  68 used  3 times (syndrom bits 42 45 52)
//  input bit  69 used  3 times (syndrom bits 49 50 53)
//  input bit  70 used  3 times (syndrom bits 36 39 46)
//  input bit  71 used  3 times (syndrom bits 43 44 47)
//  input bit  72 used  3 times (syndrom bits 30 33 40)
//  input bit  73 used  3 times (syndrom bits 37 38 41)
//  input bit  74 used  3 times (syndrom bits 24 27 34)
//  input bit  75 used  3 times (syndrom bits 31 32 35)
//  input bit  76 used  3 times (syndrom bits 18 21 28)
//  input bit  77 used  3 times (syndrom bits 25 26 29)
//  input bit  78 used  3 times (syndrom bits 12 15 22)
//  input bit  79 used  3 times (syndrom bits 19 20 23)
//  input bit  80 used  3 times (syndrom bits 6 9 16)
//  input bit  81 used  3 times (syndrom bits 13 14 17)
//  input bit  82 used  3 times (syndrom bits 0 3 11)
//  input bit  83 used  3 times (syndrom bits 7 8 11)
//  input bit  84 used  3 times (syndrom bits 1 2 11)
//  input bit  85 used  3 times (syndrom bits 1 4 5)
//  input bit  86 used  3 times (syndrom bits 2 4 5)
//  input bit  87 used  3 times (syndrom bits 7 8 10)
//  input bit  88 used  3 times (syndrom bits 0 3 17)
//  input bit  89 used  3 times (syndrom bits 13 14 16)
//  input bit  90 used  3 times (syndrom bits 6 9 23)
//  input bit  91 used  3 times (syndrom bits 19 20 22)
//  input bit  92 used  3 times (syndrom bits 12 15 29)
//  input bit  93 used  3 times (syndrom bits 25 26 28)
//  input bit  94 used  3 times (syndrom bits 18 21 35)
//  input bit  95 used  3 times (syndrom bits 31 32 34)
//  input bit  96 used  3 times (syndrom bits 24 27 41)
//  input bit  97 used  3 times (syndrom bits 37 38 40)
//  input bit  98 used  3 times (syndrom bits 30 33 47)
//  input bit  99 used  3 times (syndrom bits 43 44 46)
//  input bit 100 used  3 times (syndrom bits 36 39 53)
//  input bit 101 used  3 times (syndrom bits 49 50 52)
//  input bit 102 used  3 times (syndrom bits 42 45 59)
//  input bit 103 used  3 times (syndrom bits 55 56 58)
//  input bit 104 used  3 times (syndrom bits 48 51 61)
//  input bit 105 used  3 times (syndrom bits 60 62 63)
//  input bit 106 used  3 times (syndrom bits 54 57 63)
//  input bit 107 used  3 times (syndrom bits 54 57 62)
//  input bit 108 used  3 times (syndrom bits 48 51 60)
//  input bit 109 used  3 times (syndrom bits 55 56 61)
//  input bit 110 used  3 times (syndrom bits 42 45 58)
//  input bit 111 used  3 times (syndrom bits 49 50 59)
//  input bit 112 used  3 times (syndrom bits 36 39 52)
//  input bit 113 used  3 times (syndrom bits 43 44 53)
//  input bit 114 used  3 times (syndrom bits 30 33 46)
//  input bit 115 used  3 times (syndrom bits 37 38 47)
//  input bit 116 used  3 times (syndrom bits 24 27 40)
//  input bit 117 used  3 times (syndrom bits 31 32 41)
//  input bit 118 used  3 times (syndrom bits 18 21 34)
//  input bit 119 used  3 times (syndrom bits 25 26 35)
//  input bit 120 used  3 times (syndrom bits 12 15 28)
//  input bit 121 used  3 times (syndrom bits 19 20 29)
//  input bit 122 used  3 times (syndrom bits 6 9 22)
//  input bit 123 used  3 times (syndrom bits 13 14 23)
//  input bit 124 used  3 times (syndrom bits 0 3 16)
//  input bit 125 used  3 times (syndrom bits 7 8 17)
//  input bit 126 used  3 times (syndrom bits 4 5 10)
//  input bit 127 used  3 times (syndrom bits 1 2 10)
function [64-1:0] extended_hamming_code_192_128_f;
    input [128-1:0] in;
    reg [64-1:0] syndrom;
    begin
        syndrom[ 0] = in[  0]^in[ 41]^in[ 44]^in[ 82]^in[ 88]^in[124];//6 inputs
        syndrom[ 1] = in[  0]^in[ 42]^in[ 43]^in[ 84]^in[ 85]^in[127];//6 inputs
        syndrom[ 2] = in[  0]^in[ 42]^in[ 43]^in[ 84]^in[ 86]^in[127];//6 inputs
        syndrom[ 3] = in[  1]^in[ 40]^in[ 45]^in[ 82]^in[ 88]^in[124];//6 inputs
        syndrom[ 4] = in[  1]^in[ 41]^in[ 42]^in[ 85]^in[ 86]^in[126];//6 inputs
        syndrom[ 5] = in[  1]^in[ 41]^in[ 43]^in[ 85]^in[ 86]^in[126];//6 inputs
        syndrom[ 6] = in[  2]^in[ 39]^in[ 46]^in[ 80]^in[ 90]^in[122];//6 inputs
        syndrom[ 7] = in[  2]^in[ 40]^in[ 44]^in[ 83]^in[ 87]^in[125];//6 inputs
        syndrom[ 8] = in[  2]^in[ 40]^in[ 44]^in[ 83]^in[ 87]^in[125];//6 inputs
        syndrom[ 9] = in[  3]^in[ 38]^in[ 47]^in[ 80]^in[ 90]^in[122];//6 inputs
        syndrom[10] = in[  3]^in[ 39]^in[ 45]^in[ 87]^in[126]^in[127];//6 inputs
        syndrom[11] = in[  3]^in[ 39]^in[ 45]^in[ 82]^in[ 83]^in[ 84];//6 inputs
        syndrom[12] = in[  4]^in[ 37]^in[ 48]^in[ 78]^in[ 92]^in[120];//6 inputs
        syndrom[13] = in[  4]^in[ 38]^in[ 46]^in[ 81]^in[ 89]^in[123];//6 inputs
        syndrom[14] = in[  4]^in[ 38]^in[ 46]^in[ 81]^in[ 89]^in[123];//6 inputs
        syndrom[15] = in[  5]^in[ 36]^in[ 49]^in[ 78]^in[ 92]^in[120];//6 inputs
        syndrom[16] = in[  5]^in[ 37]^in[ 47]^in[ 80]^in[ 89]^in[124];//6 inputs
        syndrom[17] = in[  5]^in[ 37]^in[ 47]^in[ 81]^in[ 88]^in[125];//6 inputs
        syndrom[18] = in[  6]^in[ 35]^in[ 50]^in[ 76]^in[ 94]^in[118];//6 inputs
        syndrom[19] = in[  6]^in[ 36]^in[ 48]^in[ 79]^in[ 91]^in[121];//6 inputs
        syndrom[20] = in[  6]^in[ 36]^in[ 48]^in[ 79]^in[ 91]^in[121];//6 inputs
        syndrom[21] = in[  7]^in[ 34]^in[ 51]^in[ 76]^in[ 94]^in[118];//6 inputs
        syndrom[22] = in[  7]^in[ 35]^in[ 49]^in[ 78]^in[ 91]^in[122];//6 inputs
        syndrom[23] = in[  7]^in[ 35]^in[ 49]^in[ 79]^in[ 90]^in[123];//6 inputs
        syndrom[24] = in[  8]^in[ 33]^in[ 52]^in[ 74]^in[ 96]^in[116];//6 inputs
        syndrom[25] = in[  8]^in[ 34]^in[ 50]^in[ 77]^in[ 93]^in[119];//6 inputs
        syndrom[26] = in[  8]^in[ 34]^in[ 50]^in[ 77]^in[ 93]^in[119];//6 inputs
        syndrom[27] = in[  9]^in[ 32]^in[ 53]^in[ 74]^in[ 96]^in[116];//6 inputs
        syndrom[28] = in[  9]^in[ 33]^in[ 51]^in[ 76]^in[ 93]^in[120];//6 inputs
        syndrom[29] = in[  9]^in[ 33]^in[ 51]^in[ 77]^in[ 92]^in[121];//6 inputs
        syndrom[30] = in[ 10]^in[ 31]^in[ 54]^in[ 72]^in[ 98]^in[114];//6 inputs
        syndrom[31] = in[ 10]^in[ 32]^in[ 52]^in[ 75]^in[ 95]^in[117];//6 inputs
        syndrom[32] = in[ 10]^in[ 32]^in[ 52]^in[ 75]^in[ 95]^in[117];//6 inputs
        syndrom[33] = in[ 11]^in[ 30]^in[ 55]^in[ 72]^in[ 98]^in[114];//6 inputs
        syndrom[34] = in[ 11]^in[ 31]^in[ 53]^in[ 74]^in[ 95]^in[118];//6 inputs
        syndrom[35] = in[ 11]^in[ 31]^in[ 53]^in[ 75]^in[ 94]^in[119];//6 inputs
        syndrom[36] = in[ 12]^in[ 29]^in[ 56]^in[ 70]^in[100]^in[112];//6 inputs
        syndrom[37] = in[ 12]^in[ 30]^in[ 54]^in[ 73]^in[ 97]^in[115];//6 inputs
        syndrom[38] = in[ 12]^in[ 30]^in[ 54]^in[ 73]^in[ 97]^in[115];//6 inputs
        syndrom[39] = in[ 13]^in[ 28]^in[ 57]^in[ 70]^in[100]^in[112];//6 inputs
        syndrom[40] = in[ 13]^in[ 29]^in[ 55]^in[ 72]^in[ 97]^in[116];//6 inputs
        syndrom[41] = in[ 13]^in[ 29]^in[ 55]^in[ 73]^in[ 96]^in[117];//6 inputs
        syndrom[42] = in[ 14]^in[ 27]^in[ 58]^in[ 68]^in[102]^in[110];//6 inputs
        syndrom[43] = in[ 14]^in[ 28]^in[ 56]^in[ 71]^in[ 99]^in[113];//6 inputs
        syndrom[44] = in[ 14]^in[ 28]^in[ 56]^in[ 71]^in[ 99]^in[113];//6 inputs
        syndrom[45] = in[ 15]^in[ 26]^in[ 59]^in[ 68]^in[102]^in[110];//6 inputs
        syndrom[46] = in[ 15]^in[ 27]^in[ 57]^in[ 70]^in[ 99]^in[114];//6 inputs
        syndrom[47] = in[ 15]^in[ 27]^in[ 57]^in[ 71]^in[ 98]^in[115];//6 inputs
        syndrom[48] = in[ 16]^in[ 25]^in[ 60]^in[ 66]^in[104]^in[108];//6 inputs
        syndrom[49] = in[ 16]^in[ 26]^in[ 58]^in[ 69]^in[101]^in[111];//6 inputs
        syndrom[50] = in[ 16]^in[ 26]^in[ 58]^in[ 69]^in[101]^in[111];//6 inputs
        syndrom[51] = in[ 17]^in[ 24]^in[ 61]^in[ 66]^in[104]^in[108];//6 inputs
        syndrom[52] = in[ 17]^in[ 25]^in[ 59]^in[ 68]^in[101]^in[112];//6 inputs
        syndrom[53] = in[ 17]^in[ 25]^in[ 59]^in[ 69]^in[100]^in[113];//6 inputs
        syndrom[54] = in[ 18]^in[ 23]^in[ 62]^in[ 64]^in[106]^in[107];//6 inputs
        syndrom[55] = in[ 18]^in[ 24]^in[ 60]^in[ 67]^in[103]^in[109];//6 inputs
        syndrom[56] = in[ 18]^in[ 24]^in[ 60]^in[ 67]^in[103]^in[109];//6 inputs
        syndrom[57] = in[ 19]^in[ 22]^in[ 63]^in[ 64]^in[106]^in[107];//6 inputs
        syndrom[58] = in[ 19]^in[ 23]^in[ 61]^in[ 66]^in[103]^in[110];//6 inputs
        syndrom[59] = in[ 19]^in[ 23]^in[ 61]^in[ 67]^in[102]^in[111];//6 inputs
        syndrom[60] = in[ 20]^in[ 21]^in[ 63]^in[ 64]^in[105]^in[108];//6 inputs
        syndrom[61] = in[ 20]^in[ 21]^in[ 63]^in[ 65]^in[104]^in[109];//6 inputs
        syndrom[62] = in[ 20]^in[ 22]^in[ 62]^in[ 65]^in[105]^in[107];//6 inputs
        syndrom[63] = in[ 21]^in[ 22]^in[ 62]^in[ 65]^in[105]^in[106];//6 inputs
        extended_hamming_code_192_128_f = syndrom;
    end
endfunction
wire [64-1:0] stored_data_edc = extended_hamming_code_192_128_f(i_stored_data);
wire [64-1:0] syndroms = i_stored_edc ^ stored_data_edc;
always @* o_detection = |syndroms;
endmodule
module ecc_ehc_128_balanced (
	input wire [128-1:0] i_write_data, // Data to write to storage
	output reg [64-1:0] o_write_edc, // EDC bits to write to storage
	input wire [128-1:0] i_stored_data, // Data read from storage, may contain error(s)
	input wire [64-1:0] i_stored_edc, // EDC bits read from storage, may conatin error(s)
	output reg [128-1:0] o_read_data, // Error free read data (as long as error was correctable)
	output reg o_correction, //indication that an error is corrected
	output reg o_detection //indication that an error is detected, this happens only if the error is not correctable
);
//extended_hamming_code_192_128_f
//Compute 64 bits Error Detection Code from a 128 bits input.
//The EDC is an extended hamming code capable of detecting any 1,2 and 3 bits errors in the input data or the EDC.
//Input usage report:
//  input bit   0 used  3 times (syndrom bits 0 1 2)
//  input bit   1 used  3 times (syndrom bits 3 4 5)
//  input bit   2 used  3 times (syndrom bits 6 7 8)
//  input bit   3 used  3 times (syndrom bits 9 10 11)
//  input bit   4 used  3 times (syndrom bits 12 13 14)
//  input bit   5 used  3 times (syndrom bits 15 16 17)
//  input bit   6 used  3 times (syndrom bits 18 19 20)
//  input bit   7 used  3 times (syndrom bits 21 22 23)
//  input bit   8 used  3 times (syndrom bits 24 25 26)
//  input bit   9 used  3 times (syndrom bits 27 28 29)
//  input bit  10 used  3 times (syndrom bits 30 31 32)
//  input bit  11 used  3 times (syndrom bits 33 34 35)
//  input bit  12 used  3 times (syndrom bits 36 37 38)
//  input bit  13 used  3 times (syndrom bits 39 40 41)
//  input bit  14 used  3 times (syndrom bits 42 43 44)
//  input bit  15 used  3 times (syndrom bits 45 46 47)
//  input bit  16 used  3 times (syndrom bits 48 49 50)
//  input bit  17 used  3 times (syndrom bits 51 52 53)
//  input bit  18 used  3 times (syndrom bits 54 55 56)
//  input bit  19 used  3 times (syndrom bits 57 58 59)
//  input bit  20 used  3 times (syndrom bits 60 61 62)
//  input bit  21 used  3 times (syndrom bits 60 61 63)
//  input bit  22 used  3 times (syndrom bits 57 62 63)
//  input bit  23 used  3 times (syndrom bits 54 58 59)
//  input bit  24 used  3 times (syndrom bits 51 55 56)
//  input bit  25 used  3 times (syndrom bits 48 52 53)
//  input bit  26 used  3 times (syndrom bits 45 49 50)
//  input bit  27 used  3 times (syndrom bits 42 46 47)
//  input bit  28 used  3 times (syndrom bits 39 43 44)
//  input bit  29 used  3 times (syndrom bits 36 40 41)
//  input bit  30 used  3 times (syndrom bits 33 37 38)
//  input bit  31 used  3 times (syndrom bits 30 34 35)
//  input bit  32 used  3 times (syndrom bits 27 31 32)
//  input bit  33 used  3 times (syndrom bits 24 28 29)
//  input bit  34 used  3 times (syndrom bits 21 25 26)
//  input bit  35 used  3 times (syndrom bits 18 22 23)
//  input bit  36 used  3 times (syndrom bits 15 19 20)
//  input bit  37 used  3 times (syndrom bits 12 16 17)
//  input bit  38 used  3 times (syndrom bits 9 13 14)
//  input bit  39 used  3 times (syndrom bits 6 10 11)
//  input bit  40 used  3 times (syndrom bits 3 7 8)
//  input bit  41 used  3 times (syndrom bits 0 4 5)
//  input bit  42 used  3 times (syndrom bits 1 2 4)
//  input bit  43 used  3 times (syndrom bits 1 2 5)
//  input bit  44 used  3 times (syndrom bits 0 7 8)
//  input bit  45 used  3 times (syndrom bits 3 10 11)
//  input bit  46 used  3 times (syndrom bits 6 13 14)
//  input bit  47 used  3 times (syndrom bits 9 16 17)
//  input bit  48 used  3 times (syndrom bits 12 19 20)
//  input bit  49 used  3 times (syndrom bits 15 22 23)
//  input bit  50 used  3 times (syndrom bits 18 25 26)
//  input bit  51 used  3 times (syndrom bits 21 28 29)
//  input bit  52 used  3 times (syndrom bits 24 31 32)
//  input bit  53 used  3 times (syndrom bits 27 34 35)
//  input bit  54 used  3 times (syndrom bits 30 37 38)
//  input bit  55 used  3 times (syndrom bits 33 40 41)
//  input bit  56 used  3 times (syndrom bits 36 43 44)
//  input bit  57 used  3 times (syndrom bits 39 46 47)
//  input bit  58 used  3 times (syndrom bits 42 49 50)
//  input bit  59 used  3 times (syndrom bits 45 52 53)
//  input bit  60 used  3 times (syndrom bits 48 55 56)
//  input bit  61 used  3 times (syndrom bits 51 58 59)
//  input bit  62 used  3 times (syndrom bits 54 62 63)
//  input bit  63 used  3 times (syndrom bits 57 60 61)
//  input bit  64 used  3 times (syndrom bits 54 57 60)
//  input bit  65 used  3 times (syndrom bits 61 62 63)
//  input bit  66 used  3 times (syndrom bits 48 51 58)
//  input bit  67 used  3 times (syndrom bits 55 56 59)
//  input bit  68 used  3 times (syndrom bits 42 45 52)
//  input bit  69 used  3 times (syndrom bits 49 50 53)
//  input bit  70 used  3 times (syndrom bits 36 39 46)
//  input bit  71 used  3 times (syndrom bits 43 44 47)
//  input bit  72 used  3 times (syndrom bits 30 33 40)
//  input bit  73 used  3 times (syndrom bits 37 38 41)
//  input bit  74 used  3 times (syndrom bits 24 27 34)
//  input bit  75 used  3 times (syndrom bits 31 32 35)
//  input bit  76 used  3 times (syndrom bits 18 21 28)
//  input bit  77 used  3 times (syndrom bits 25 26 29)
//  input bit  78 used  3 times (syndrom bits 12 15 22)
//  input bit  79 used  3 times (syndrom bits 19 20 23)
//  input bit  80 used  3 times (syndrom bits 6 9 16)
//  input bit  81 used  3 times (syndrom bits 13 14 17)
//  input bit  82 used  3 times (syndrom bits 0 3 11)
//  input bit  83 used  3 times (syndrom bits 7 8 11)
//  input bit  84 used  3 times (syndrom bits 1 2 11)
//  input bit  85 used  3 times (syndrom bits 1 4 5)
//  input bit  86 used  3 times (syndrom bits 2 4 5)
//  input bit  87 used  3 times (syndrom bits 7 8 10)
//  input bit  88 used  3 times (syndrom bits 0 3 17)
//  input bit  89 used  3 times (syndrom bits 13 14 16)
//  input bit  90 used  3 times (syndrom bits 6 9 23)
//  input bit  91 used  3 times (syndrom bits 19 20 22)
//  input bit  92 used  3 times (syndrom bits 12 15 29)
//  input bit  93 used  3 times (syndrom bits 25 26 28)
//  input bit  94 used  3 times (syndrom bits 18 21 35)
//  input bit  95 used  3 times (syndrom bits 31 32 34)
//  input bit  96 used  3 times (syndrom bits 24 27 41)
//  input bit  97 used  3 times (syndrom bits 37 38 40)
//  input bit  98 used  3 times (syndrom bits 30 33 47)
//  input bit  99 used  3 times (syndrom bits 43 44 46)
//  input bit 100 used  3 times (syndrom bits 36 39 53)
//  input bit 101 used  3 times (syndrom bits 49 50 52)
//  input bit 102 used  3 times (syndrom bits 42 45 59)
//  input bit 103 used  3 times (syndrom bits 55 56 58)
//  input bit 104 used  3 times (syndrom bits 48 51 61)
//  input bit 105 used  3 times (syndrom bits 60 62 63)
//  input bit 106 used  3 times (syndrom bits 54 57 63)
//  input bit 107 used  3 times (syndrom bits 54 57 62)
//  input bit 108 used  3 times (syndrom bits 48 51 60)
//  input bit 109 used  3 times (syndrom bits 55 56 61)
//  input bit 110 used  3 times (syndrom bits 42 45 58)
//  input bit 111 used  3 times (syndrom bits 49 50 59)
//  input bit 112 used  3 times (syndrom bits 36 39 52)
//  input bit 113 used  3 times (syndrom bits 43 44 53)
//  input bit 114 used  3 times (syndrom bits 30 33 46)
//  input bit 115 used  3 times (syndrom bits 37 38 47)
//  input bit 116 used  3 times (syndrom bits 24 27 40)
//  input bit 117 used  3 times (syndrom bits 31 32 41)
//  input bit 118 used  3 times (syndrom bits 18 21 34)
//  input bit 119 used  3 times (syndrom bits 25 26 35)
//  input bit 120 used  3 times (syndrom bits 12 15 28)
//  input bit 121 used  3 times (syndrom bits 19 20 29)
//  input bit 122 used  3 times (syndrom bits 6 9 22)
//  input bit 123 used  3 times (syndrom bits 13 14 23)
//  input bit 124 used  3 times (syndrom bits 0 3 16)
//  input bit 125 used  3 times (syndrom bits 7 8 17)
//  input bit 126 used  3 times (syndrom bits 4 5 10)
//  input bit 127 used  3 times (syndrom bits 1 2 10)
function [64-1:0] extended_hamming_code_192_128_f;
    input [128-1:0] in;
    reg [64-1:0] syndrom;
    begin
        syndrom[ 0] = in[  0]^in[ 41]^in[ 44]^in[ 82]^in[ 88]^in[124];//6 inputs
        syndrom[ 1] = in[  0]^in[ 42]^in[ 43]^in[ 84]^in[ 85]^in[127];//6 inputs
        syndrom[ 2] = in[  0]^in[ 42]^in[ 43]^in[ 84]^in[ 86]^in[127];//6 inputs
        syndrom[ 3] = in[  1]^in[ 40]^in[ 45]^in[ 82]^in[ 88]^in[124];//6 inputs
        syndrom[ 4] = in[  1]^in[ 41]^in[ 42]^in[ 85]^in[ 86]^in[126];//6 inputs
        syndrom[ 5] = in[  1]^in[ 41]^in[ 43]^in[ 85]^in[ 86]^in[126];//6 inputs
        syndrom[ 6] = in[  2]^in[ 39]^in[ 46]^in[ 80]^in[ 90]^in[122];//6 inputs
        syndrom[ 7] = in[  2]^in[ 40]^in[ 44]^in[ 83]^in[ 87]^in[125];//6 inputs
        syndrom[ 8] = in[  2]^in[ 40]^in[ 44]^in[ 83]^in[ 87]^in[125];//6 inputs
        syndrom[ 9] = in[  3]^in[ 38]^in[ 47]^in[ 80]^in[ 90]^in[122];//6 inputs
        syndrom[10] = in[  3]^in[ 39]^in[ 45]^in[ 87]^in[126]^in[127];//6 inputs
        syndrom[11] = in[  3]^in[ 39]^in[ 45]^in[ 82]^in[ 83]^in[ 84];//6 inputs
        syndrom[12] = in[  4]^in[ 37]^in[ 48]^in[ 78]^in[ 92]^in[120];//6 inputs
        syndrom[13] = in[  4]^in[ 38]^in[ 46]^in[ 81]^in[ 89]^in[123];//6 inputs
        syndrom[14] = in[  4]^in[ 38]^in[ 46]^in[ 81]^in[ 89]^in[123];//6 inputs
        syndrom[15] = in[  5]^in[ 36]^in[ 49]^in[ 78]^in[ 92]^in[120];//6 inputs
        syndrom[16] = in[  5]^in[ 37]^in[ 47]^in[ 80]^in[ 89]^in[124];//6 inputs
        syndrom[17] = in[  5]^in[ 37]^in[ 47]^in[ 81]^in[ 88]^in[125];//6 inputs
        syndrom[18] = in[  6]^in[ 35]^in[ 50]^in[ 76]^in[ 94]^in[118];//6 inputs
        syndrom[19] = in[  6]^in[ 36]^in[ 48]^in[ 79]^in[ 91]^in[121];//6 inputs
        syndrom[20] = in[  6]^in[ 36]^in[ 48]^in[ 79]^in[ 91]^in[121];//6 inputs
        syndrom[21] = in[  7]^in[ 34]^in[ 51]^in[ 76]^in[ 94]^in[118];//6 inputs
        syndrom[22] = in[  7]^in[ 35]^in[ 49]^in[ 78]^in[ 91]^in[122];//6 inputs
        syndrom[23] = in[  7]^in[ 35]^in[ 49]^in[ 79]^in[ 90]^in[123];//6 inputs
        syndrom[24] = in[  8]^in[ 33]^in[ 52]^in[ 74]^in[ 96]^in[116];//6 inputs
        syndrom[25] = in[  8]^in[ 34]^in[ 50]^in[ 77]^in[ 93]^in[119];//6 inputs
        syndrom[26] = in[  8]^in[ 34]^in[ 50]^in[ 77]^in[ 93]^in[119];//6 inputs
        syndrom[27] = in[  9]^in[ 32]^in[ 53]^in[ 74]^in[ 96]^in[116];//6 inputs
        syndrom[28] = in[  9]^in[ 33]^in[ 51]^in[ 76]^in[ 93]^in[120];//6 inputs
        syndrom[29] = in[  9]^in[ 33]^in[ 51]^in[ 77]^in[ 92]^in[121];//6 inputs
        syndrom[30] = in[ 10]^in[ 31]^in[ 54]^in[ 72]^in[ 98]^in[114];//6 inputs
        syndrom[31] = in[ 10]^in[ 32]^in[ 52]^in[ 75]^in[ 95]^in[117];//6 inputs
        syndrom[32] = in[ 10]^in[ 32]^in[ 52]^in[ 75]^in[ 95]^in[117];//6 inputs
        syndrom[33] = in[ 11]^in[ 30]^in[ 55]^in[ 72]^in[ 98]^in[114];//6 inputs
        syndrom[34] = in[ 11]^in[ 31]^in[ 53]^in[ 74]^in[ 95]^in[118];//6 inputs
        syndrom[35] = in[ 11]^in[ 31]^in[ 53]^in[ 75]^in[ 94]^in[119];//6 inputs
        syndrom[36] = in[ 12]^in[ 29]^in[ 56]^in[ 70]^in[100]^in[112];//6 inputs
        syndrom[37] = in[ 12]^in[ 30]^in[ 54]^in[ 73]^in[ 97]^in[115];//6 inputs
        syndrom[38] = in[ 12]^in[ 30]^in[ 54]^in[ 73]^in[ 97]^in[115];//6 inputs
        syndrom[39] = in[ 13]^in[ 28]^in[ 57]^in[ 70]^in[100]^in[112];//6 inputs
        syndrom[40] = in[ 13]^in[ 29]^in[ 55]^in[ 72]^in[ 97]^in[116];//6 inputs
        syndrom[41] = in[ 13]^in[ 29]^in[ 55]^in[ 73]^in[ 96]^in[117];//6 inputs
        syndrom[42] = in[ 14]^in[ 27]^in[ 58]^in[ 68]^in[102]^in[110];//6 inputs
        syndrom[43] = in[ 14]^in[ 28]^in[ 56]^in[ 71]^in[ 99]^in[113];//6 inputs
        syndrom[44] = in[ 14]^in[ 28]^in[ 56]^in[ 71]^in[ 99]^in[113];//6 inputs
        syndrom[45] = in[ 15]^in[ 26]^in[ 59]^in[ 68]^in[102]^in[110];//6 inputs
        syndrom[46] = in[ 15]^in[ 27]^in[ 57]^in[ 70]^in[ 99]^in[114];//6 inputs
        syndrom[47] = in[ 15]^in[ 27]^in[ 57]^in[ 71]^in[ 98]^in[115];//6 inputs
        syndrom[48] = in[ 16]^in[ 25]^in[ 60]^in[ 66]^in[104]^in[108];//6 inputs
        syndrom[49] = in[ 16]^in[ 26]^in[ 58]^in[ 69]^in[101]^in[111];//6 inputs
        syndrom[50] = in[ 16]^in[ 26]^in[ 58]^in[ 69]^in[101]^in[111];//6 inputs
        syndrom[51] = in[ 17]^in[ 24]^in[ 61]^in[ 66]^in[104]^in[108];//6 inputs
        syndrom[52] = in[ 17]^in[ 25]^in[ 59]^in[ 68]^in[101]^in[112];//6 inputs
        syndrom[53] = in[ 17]^in[ 25]^in[ 59]^in[ 69]^in[100]^in[113];//6 inputs
        syndrom[54] = in[ 18]^in[ 23]^in[ 62]^in[ 64]^in[106]^in[107];//6 inputs
        syndrom[55] = in[ 18]^in[ 24]^in[ 60]^in[ 67]^in[103]^in[109];//6 inputs
        syndrom[56] = in[ 18]^in[ 24]^in[ 60]^in[ 67]^in[103]^in[109];//6 inputs
        syndrom[57] = in[ 19]^in[ 22]^in[ 63]^in[ 64]^in[106]^in[107];//6 inputs
        syndrom[58] = in[ 19]^in[ 23]^in[ 61]^in[ 66]^in[103]^in[110];//6 inputs
        syndrom[59] = in[ 19]^in[ 23]^in[ 61]^in[ 67]^in[102]^in[111];//6 inputs
        syndrom[60] = in[ 20]^in[ 21]^in[ 63]^in[ 64]^in[105]^in[108];//6 inputs
        syndrom[61] = in[ 20]^in[ 21]^in[ 63]^in[ 65]^in[104]^in[109];//6 inputs
        syndrom[62] = in[ 20]^in[ 22]^in[ 62]^in[ 65]^in[105]^in[107];//6 inputs
        syndrom[63] = in[ 21]^in[ 22]^in[ 62]^in[ 65]^in[105]^in[106];//6 inputs
        extended_hamming_code_192_128_f = syndrom;
    end
endfunction
function [2+128-1:0] extended_hamming_code_192_128_f_correction_pattern_f;
    input [64-1:0] syndrom;
	input correctEdcSingleBitErrors;
	reg uncorrectable_error;
	reg correctable_error;
	reg [128-1:0] correction_pattern;
	reg edcSingleBitErrorFillValue;
    begin
		edcSingleBitErrorFillValue = correctEdcSingleBitErrors ? 1'b0 : 1'bx;
		correction_pattern = {128{1'bx}};
		correctable_error = 1'b1;
        uncorrectable_error = 1'b0;
		case(syndrom)
			64'b0000000000000000000000000000000000000000000000000000000000000000: begin
				correctable_error = 1'b0;
				correction_pattern = {128{1'b0}};
			end	
			64'b0000000000000000000000000000000000000000000000000000000000000111: begin
				correction_pattern = {128{1'b0}};correction_pattern[  0]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000111000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  1]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000111000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  2]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000111000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  3]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000111000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  4]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000111000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  5]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000111000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  6]=1'b1;
			end
			64'b0000000000000000000000000000000000000000111000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  7]=1'b1;
			end
			64'b0000000000000000000000000000000000000111000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  8]=1'b1;
			end
			64'b0000000000000000000000000000000000111000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[  9]=1'b1;
			end
			64'b0000000000000000000000000000000111000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 10]=1'b1;
			end
			64'b0000000000000000000000000000111000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 11]=1'b1;
			end
			64'b0000000000000000000000000111000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 12]=1'b1;
			end
			64'b0000000000000000000000111000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 13]=1'b1;
			end
			64'b0000000000000000000111000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 14]=1'b1;
			end
			64'b0000000000000000111000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 15]=1'b1;
			end
			64'b0000000000000111000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 16]=1'b1;
			end
			64'b0000000000111000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 17]=1'b1;
			end
			64'b0000000111000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 18]=1'b1;
			end
			64'b0000111000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 19]=1'b1;
			end
			64'b0111000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 20]=1'b1;
			end
			64'b1011000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 21]=1'b1;
			end
			64'b1100001000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 22]=1'b1;
			end
			64'b0000110001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 23]=1'b1;
			end
			64'b0000000110001000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 24]=1'b1;
			end
			64'b0000000000110001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 25]=1'b1;
			end
			64'b0000000000000110001000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 26]=1'b1;
			end
			64'b0000000000000000110001000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 27]=1'b1;
			end
			64'b0000000000000000000110001000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 28]=1'b1;
			end
			64'b0000000000000000000000110001000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 29]=1'b1;
			end
			64'b0000000000000000000000000110001000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 30]=1'b1;
			end
			64'b0000000000000000000000000000110001000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 31]=1'b1;
			end
			64'b0000000000000000000000000000000110001000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 32]=1'b1;
			end
			64'b0000000000000000000000000000000000110001000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 33]=1'b1;
			end
			64'b0000000000000000000000000000000000000110001000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 34]=1'b1;
			end
			64'b0000000000000000000000000000000000000000110001000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 35]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000110001000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 36]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000110001000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 37]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000110001000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 38]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000110001000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 39]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000110001000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 40]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000110001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 41]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000010110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 42]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000100110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 43]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000110000001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 44]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000110000001000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 45]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000110000001000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 46]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000110000001000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 47]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000110000001000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 48]=1'b1;
			end
			64'b0000000000000000000000000000000000000000110000001000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 49]=1'b1;
			end
			64'b0000000000000000000000000000000000000110000001000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 50]=1'b1;
			end
			64'b0000000000000000000000000000000000110000001000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 51]=1'b1;
			end
			64'b0000000000000000000000000000000110000001000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 52]=1'b1;
			end
			64'b0000000000000000000000000000110000001000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 53]=1'b1;
			end
			64'b0000000000000000000000000110000001000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 54]=1'b1;
			end
			64'b0000000000000000000000110000001000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 55]=1'b1;
			end
			64'b0000000000000000000110000001000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 56]=1'b1;
			end
			64'b0000000000000000110000001000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 57]=1'b1;
			end
			64'b0000000000000110000001000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 58]=1'b1;
			end
			64'b0000000000110000001000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 59]=1'b1;
			end
			64'b0000000110000001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 60]=1'b1;
			end
			64'b0000110000001000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 61]=1'b1;
			end
			64'b1100000001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 62]=1'b1;
			end
			64'b0011001000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 63]=1'b1;
			end
			64'b0001001001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 64]=1'b1;
			end
			64'b1110000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 65]=1'b1;
			end
			64'b0000010000001001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 66]=1'b1;
			end
			64'b0000100110000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 67]=1'b1;
			end
			64'b0000000000010000001001000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 68]=1'b1;
			end
			64'b0000000000100110000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 69]=1'b1;
			end
			64'b0000000000000000010000001001000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 70]=1'b1;
			end
			64'b0000000000000000100110000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 71]=1'b1;
			end
			64'b0000000000000000000000010000001001000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 72]=1'b1;
			end
			64'b0000000000000000000000100110000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 73]=1'b1;
			end
			64'b0000000000000000000000000000010000001001000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 74]=1'b1;
			end
			64'b0000000000000000000000000000100110000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 75]=1'b1;
			end
			64'b0000000000000000000000000000000000010000001001000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 76]=1'b1;
			end
			64'b0000000000000000000000000000000000100110000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 77]=1'b1;
			end
			64'b0000000000000000000000000000000000000000010000001001000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 78]=1'b1;
			end
			64'b0000000000000000000000000000000000000000100110000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 79]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000010000001001000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 80]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000100110000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 81]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000100000001001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 82]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000100110000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 83]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000100000000110: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 84]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000110010: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 85]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000110100: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 86]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000010110000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 87]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000100000000000001001: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 88]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000010110000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 89]=1'b1;
			end
			64'b0000000000000000000000000000000000000000100000000000001001000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 90]=1'b1;
			end
			64'b0000000000000000000000000000000000000000010110000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 91]=1'b1;
			end
			64'b0000000000000000000000000000000000100000000000001001000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 92]=1'b1;
			end
			64'b0000000000000000000000000000000000010110000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 93]=1'b1;
			end
			64'b0000000000000000000000000000100000000000001001000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 94]=1'b1;
			end
			64'b0000000000000000000000000000010110000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 95]=1'b1;
			end
			64'b0000000000000000000000100000000000001001000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 96]=1'b1;
			end
			64'b0000000000000000000000010110000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 97]=1'b1;
			end
			64'b0000000000000000100000000000001001000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 98]=1'b1;
			end
			64'b0000000000000000010110000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[ 99]=1'b1;
			end
			64'b0000000000100000000000001001000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[100]=1'b1;
			end
			64'b0000000000010110000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[101]=1'b1;
			end
			64'b0000100000000000001001000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[102]=1'b1;
			end
			64'b0000010110000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[103]=1'b1;
			end
			64'b0010000000001001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[104]=1'b1;
			end
			64'b1101000000000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[105]=1'b1;
			end
			64'b1000001001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[106]=1'b1;
			end
			64'b0100001001000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[107]=1'b1;
			end
			64'b0001000000001001000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[108]=1'b1;
			end
			64'b0010000110000000000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[109]=1'b1;
			end
			64'b0000010000000000001001000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[110]=1'b1;
			end
			64'b0000100000000110000000000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[111]=1'b1;
			end
			64'b0000000000010000000000001001000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[112]=1'b1;
			end
			64'b0000000000100000000110000000000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[113]=1'b1;
			end
			64'b0000000000000000010000000000001001000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[114]=1'b1;
			end
			64'b0000000000000000100000000110000000000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[115]=1'b1;
			end
			64'b0000000000000000000000010000000000001001000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[116]=1'b1;
			end
			64'b0000000000000000000000100000000110000000000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[117]=1'b1;
			end
			64'b0000000000000000000000000000010000000000001001000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[118]=1'b1;
			end
			64'b0000000000000000000000000000100000000110000000000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[119]=1'b1;
			end
			64'b0000000000000000000000000000000000010000000000001001000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[120]=1'b1;
			end
			64'b0000000000000000000000000000000000100000000110000000000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[121]=1'b1;
			end
			64'b0000000000000000000000000000000000000000010000000000001001000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[122]=1'b1;
			end
			64'b0000000000000000000000000000000000000000100000000110000000000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[123]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000010000000000001001: begin
				correction_pattern = {128{1'b0}};correction_pattern[124]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000100000000110000000: begin
				correction_pattern = {128{1'b0}};correction_pattern[125]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000010000110000: begin
				correction_pattern = {128{1'b0}};correction_pattern[126]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000010000000110: begin
				correction_pattern = {128{1'b0}};correction_pattern[127]=1'b1;
			end
			64'b0000000000000000000000000000000000000000000000000000000000000001: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000000010: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000000100: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000001000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000010000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000000100000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000001000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000010000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000000100000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000001000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000010000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000000100000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000001000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000010000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000000100000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000001000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000010000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000000100000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000001000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000010000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000000100000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000001000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000010000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000000100000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000001000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000010000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000000100000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000001000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000010000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000000100000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000001000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000010000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000000100000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000001000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000010000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000000100000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000001000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000010000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000000100000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000001000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000010000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000000100000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000001000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000010000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000000100000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000001000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000010000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000000100000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000001000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000010000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000000100000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000001000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000010000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000000100000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000001000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000010000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000000100000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000001000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000010000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0000100000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0001000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0010000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b0100000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			64'b1000000000000000000000000000000000000000000000000000000000000000: begin
				uncorrectable_error = ~correctEdcSingleBitErrors;//if we don't correct it, count it as a detected error
				correction_pattern = {128{edcSingleBitErrorFillValue}};//single bit error on EDC bits -> nothing to correct!
			end
			default: begin
				uncorrectable_error = 1'b1;
				correctable_error = 1'b0;
			end
		endcase
		extended_hamming_code_192_128_f_correction_pattern_f = {uncorrectable_error,correctable_error,correction_pattern};
    end
endfunction

wire [64-1:0] stored_data_edc = extended_hamming_code_192_128_f(i_stored_data);
wire [64-1:0] syndroms = i_stored_edc ^ stored_data_edc;
reg uncorrectable_error;
reg [128-1:0] correction_pattern;
always @* begin
	{o_detection,o_correction,correction_pattern} = extended_hamming_code_192_128_f_correction_pattern_f(syndroms,CORRECT_EDC_SINGLE_BIT_ERRORS);     
	o_read_data = i_stored_data ^ correction_pattern;
end
endmodule



